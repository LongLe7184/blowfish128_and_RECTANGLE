//R MACROS
