//-----------------------------------------------------------
// Header: Blowfish-128's Definition
//-----------------------------------------------------------
// Author	: Long Le, Manh Nguyen
// Date  	: Feb-11th, 2025
// Description	: Contain Macros holding S-Boxes's values
//-----------------------------------------------------------


//SBox1 Macro's Values
`define SBOX1_ELEMENT_000 32'hD1310BA6
`define SBOX1_ELEMENT_001 32'h98DFB5AC
`define SBOX1_ELEMENT_002 32'h2FFD72DB
`define SBOX1_ELEMENT_003 32'hD01ADFB7
`define SBOX1_ELEMENT_004 32'hB8E1AFED
`define SBOX1_ELEMENT_005 32'h6A267E96
`define SBOX1_ELEMENT_006 32'hBA7C9045
`define SBOX1_ELEMENT_007 32'hF12C7F99
`define SBOX1_ELEMENT_008 32'h24A19947
`define SBOX1_ELEMENT_009 32'hB3916CF7
`define SBOX1_ELEMENT_010 32'h0801F2E2
`define SBOX1_ELEMENT_011 32'h858EFC16
`define SBOX1_ELEMENT_012 32'h636920D8
`define SBOX1_ELEMENT_013 32'h71574E69
`define SBOX1_ELEMENT_014 32'hA458FEA3
`define SBOX1_ELEMENT_015 32'hF4933D7E
`define SBOX1_ELEMENT_016 32'h0D95748F
`define SBOX1_ELEMENT_017 32'h728EB658
`define SBOX1_ELEMENT_018 32'h718BCD58
`define SBOX1_ELEMENT_019 32'h82154AEE
`define SBOX1_ELEMENT_020 32'h7B54A41D
`define SBOX1_ELEMENT_021 32'hC25A59B5
`define SBOX1_ELEMENT_022 32'h9C30D539
`define SBOX1_ELEMENT_023 32'h2AF26013
`define SBOX1_ELEMENT_024 32'hC5D1B023
`define SBOX1_ELEMENT_025 32'h286085F0
`define SBOX1_ELEMENT_026 32'hCA417918
`define SBOX1_ELEMENT_027 32'hB8DB38EF
`define SBOX1_ELEMENT_028 32'h8E79DCB0
`define SBOX1_ELEMENT_029 32'h603A180E
`define SBOX1_ELEMENT_030 32'h6C9E0E8B
`define SBOX1_ELEMENT_031 32'hB01E8A3E
`define SBOX1_ELEMENT_032 32'hD71577C1
`define SBOX1_ELEMENT_033 32'hBD314B27
`define SBOX1_ELEMENT_034 32'h78AF2FDA
`define SBOX1_ELEMENT_035 32'h55605C60
`define SBOX1_ELEMENT_036 32'hE65525F3
`define SBOX1_ELEMENT_037 32'hAA55AB94
`define SBOX1_ELEMENT_038 32'h57489862
`define SBOX1_ELEMENT_039 32'h63E81440
`define SBOX1_ELEMENT_040 32'h55CA396A
`define SBOX1_ELEMENT_041 32'h2AAB10B6
`define SBOX1_ELEMENT_042 32'hB4CC5C34
`define SBOX1_ELEMENT_043 32'h1141E8CE
`define SBOX1_ELEMENT_044 32'hA15486AF
`define SBOX1_ELEMENT_045 32'h7C72E993
`define SBOX1_ELEMENT_046 32'hB3EE1411
`define SBOX1_ELEMENT_047 32'h636FBC2A
`define SBOX1_ELEMENT_048 32'h2BA9C55D
`define SBOX1_ELEMENT_049 32'h741831F6
`define SBOX1_ELEMENT_050 32'hCE5C3E16
`define SBOX1_ELEMENT_051 32'h9B87931E
`define SBOX1_ELEMENT_052 32'hAFD6BA33
`define SBOX1_ELEMENT_053 32'h6C24CF5C
`define SBOX1_ELEMENT_054 32'h7A325381
`define SBOX1_ELEMENT_055 32'h28958677
`define SBOX1_ELEMENT_056 32'h3B8F4898
`define SBOX1_ELEMENT_057 32'h6B4BB9AF
`define SBOX1_ELEMENT_058 32'hC4BFE81B
`define SBOX1_ELEMENT_059 32'h66282193
`define SBOX1_ELEMENT_060 32'h61D809CC
`define SBOX1_ELEMENT_061 32'hFB21A991
`define SBOX1_ELEMENT_062 32'h487CAC60
`define SBOX1_ELEMENT_063 32'h5DEC8032
`define SBOX1_ELEMENT_064 32'hEF845D5D
`define SBOX1_ELEMENT_065 32'hE98575B1
`define SBOX1_ELEMENT_066 32'hDC262302
`define SBOX1_ELEMENT_067 32'hEB651B88
`define SBOX1_ELEMENT_068 32'h23893E81
`define SBOX1_ELEMENT_069 32'hD396ACC5
`define SBOX1_ELEMENT_070 32'h0F6D6FF3
`define SBOX1_ELEMENT_071 32'h83F44239
`define SBOX1_ELEMENT_072 32'h2E0B4482
`define SBOX1_ELEMENT_073 32'hA4842004
`define SBOX1_ELEMENT_074 32'h69C8F04A
`define SBOX1_ELEMENT_075 32'h9E1F9B5E
`define SBOX1_ELEMENT_076 32'h21C66842
`define SBOX1_ELEMENT_077 32'hF6E96C9A
`define SBOX1_ELEMENT_078 32'h670C9C61
`define SBOX1_ELEMENT_079 32'hABD388F0
`define SBOX1_ELEMENT_080 32'h6A51A0D2
`define SBOX1_ELEMENT_081 32'hD8542F68
`define SBOX1_ELEMENT_082 32'h960FA728
`define SBOX1_ELEMENT_083 32'hAB5133A3
`define SBOX1_ELEMENT_084 32'h6EEF0B6C
`define SBOX1_ELEMENT_085 32'h137A3BE4
`define SBOX1_ELEMENT_086 32'hBA3BF050
`define SBOX1_ELEMENT_087 32'h7EFB2A98
`define SBOX1_ELEMENT_088 32'hA1F1651D
`define SBOX1_ELEMENT_089 32'h39AF0176
`define SBOX1_ELEMENT_090 32'h66CA593E
`define SBOX1_ELEMENT_091 32'h82430E88
`define SBOX1_ELEMENT_092 32'h8CEE8619
`define SBOX1_ELEMENT_093 32'h456F9FB4
`define SBOX1_ELEMENT_094 32'h7D84A5C3
`define SBOX1_ELEMENT_095 32'h3B8B5EBE
`define SBOX1_ELEMENT_096 32'hE06F75D8
`define SBOX1_ELEMENT_097 32'h85C12073
`define SBOX1_ELEMENT_098 32'h401A449F
`define SBOX1_ELEMENT_099 32'h56C16AA6
`define SBOX1_ELEMENT_100 32'h4ED3AA62
`define SBOX1_ELEMENT_101 32'h363F7706
`define SBOX1_ELEMENT_102 32'h1BFEDF72
`define SBOX1_ELEMENT_103 32'h429B023D
`define SBOX1_ELEMENT_104 32'h37D0D724
`define SBOX1_ELEMENT_105 32'hD00A1248
`define SBOX1_ELEMENT_106 32'hDB0FEAD3
`define SBOX1_ELEMENT_107 32'h49F1C09B
`define SBOX1_ELEMENT_108 32'h075372C9
`define SBOX1_ELEMENT_109 32'h80991B7B
`define SBOX1_ELEMENT_110 32'h25D479D8
`define SBOX1_ELEMENT_111 32'hF6E8DEF7
`define SBOX1_ELEMENT_112 32'hE3FE501A
`define SBOX1_ELEMENT_113 32'hB6794C3B
`define SBOX1_ELEMENT_114 32'h976CE0BD
`define SBOX1_ELEMENT_115 32'h04C006BA
`define SBOX1_ELEMENT_116 32'hC1A94FB6
`define SBOX1_ELEMENT_117 32'h409F60C4
`define SBOX1_ELEMENT_118 32'h5E5C9EC2
`define SBOX1_ELEMENT_119 32'h196A2463
`define SBOX1_ELEMENT_120 32'h68FB6FAF
`define SBOX1_ELEMENT_121 32'h3E6C53B5
`define SBOX1_ELEMENT_122 32'h1339B2EB
`define SBOX1_ELEMENT_123 32'h3B52EC6F
`define SBOX1_ELEMENT_124 32'h6DFC511F
`define SBOX1_ELEMENT_125 32'h9B30952C
`define SBOX1_ELEMENT_126 32'hCC814544
`define SBOX1_ELEMENT_127 32'hAF5EBD09
`define SBOX1_ELEMENT_128 32'hBEE3D004
`define SBOX1_ELEMENT_129 32'hDE334AFD
`define SBOX1_ELEMENT_130 32'h660F2807
`define SBOX1_ELEMENT_131 32'h192E4BB3
`define SBOX1_ELEMENT_132 32'hC0CBA857
`define SBOX1_ELEMENT_133 32'h45C8740F
`define SBOX1_ELEMENT_134 32'hD20B5F39
`define SBOX1_ELEMENT_135 32'hB9D3FBDB
`define SBOX1_ELEMENT_136 32'h5579C0BD
`define SBOX1_ELEMENT_137 32'h1A60320A
`define SBOX1_ELEMENT_138 32'hD6A100C6
`define SBOX1_ELEMENT_139 32'h402C7279
`define SBOX1_ELEMENT_140 32'h679F25FE
`define SBOX1_ELEMENT_141 32'hFB1FA3CC
`define SBOX1_ELEMENT_142 32'h8EA5E9F8
`define SBOX1_ELEMENT_143 32'hDB3222F8
`define SBOX1_ELEMENT_144 32'h3C7516DF
`define SBOX1_ELEMENT_145 32'hFD616B15
`define SBOX1_ELEMENT_146 32'h2F501EC8
`define SBOX1_ELEMENT_147 32'hAD0552AB
`define SBOX1_ELEMENT_148 32'h323DB5FA
`define SBOX1_ELEMENT_149 32'hFD238760
`define SBOX1_ELEMENT_150 32'h53317B48
`define SBOX1_ELEMENT_151 32'h3E00DF82
`define SBOX1_ELEMENT_152 32'h9E5C57BB
`define SBOX1_ELEMENT_153 32'hCA6F8CA0
`define SBOX1_ELEMENT_154 32'h1A87562E
`define SBOX1_ELEMENT_155 32'hDF1769DB
`define SBOX1_ELEMENT_156 32'hD542A8F6
`define SBOX1_ELEMENT_157 32'h287EFFC3
`define SBOX1_ELEMENT_158 32'hAC6732C6
`define SBOX1_ELEMENT_159 32'h8C4F5573
`define SBOX1_ELEMENT_160 32'h695B27B0
`define SBOX1_ELEMENT_161 32'hBBCA58C8
`define SBOX1_ELEMENT_162 32'hE1FFA35D
`define SBOX1_ELEMENT_163 32'hB8F011A0
`define SBOX1_ELEMENT_164 32'h10FA3D98
`define SBOX1_ELEMENT_165 32'hFD2183B8
`define SBOX1_ELEMENT_166 32'h4AFCB56C
`define SBOX1_ELEMENT_167 32'h2DD1D35B
`define SBOX1_ELEMENT_168 32'h9A53E479
`define SBOX1_ELEMENT_169 32'hB6F84565
`define SBOX1_ELEMENT_170 32'hD28E49BC
`define SBOX1_ELEMENT_171 32'h4BFB9790
`define SBOX1_ELEMENT_172 32'hE1DDF2DA
`define SBOX1_ELEMENT_173 32'hA4CB7E33
`define SBOX1_ELEMENT_174 32'h62FB1341
`define SBOX1_ELEMENT_175 32'hCEE4C6E8
`define SBOX1_ELEMENT_176 32'hEF20CADA
`define SBOX1_ELEMENT_177 32'h36774C01
`define SBOX1_ELEMENT_178 32'hD07E9EFE
`define SBOX1_ELEMENT_179 32'h2BF11FB4
`define SBOX1_ELEMENT_180 32'h95DBDA4D
`define SBOX1_ELEMENT_181 32'hAE909198
`define SBOX1_ELEMENT_182 32'hEAAD8E71
`define SBOX1_ELEMENT_183 32'h6B93D5A0
`define SBOX1_ELEMENT_184 32'hD08ED1D0
`define SBOX1_ELEMENT_185 32'hAFC725E0
`define SBOX1_ELEMENT_186 32'h8E3C5B2F
`define SBOX1_ELEMENT_187 32'h8E7594B7
`define SBOX1_ELEMENT_188 32'h8FF6E2FB
`define SBOX1_ELEMENT_189 32'hF2122B64
`define SBOX1_ELEMENT_190 32'h8888B812
`define SBOX1_ELEMENT_191 32'h900DF01C
`define SBOX1_ELEMENT_192 32'h4FAD5EA0
`define SBOX1_ELEMENT_193 32'h688FC31C
`define SBOX1_ELEMENT_194 32'hD1CFF191
`define SBOX1_ELEMENT_195 32'hB3A8C1AD
`define SBOX1_ELEMENT_196 32'h2F2F2218
`define SBOX1_ELEMENT_197 32'hBE0E1777
`define SBOX1_ELEMENT_198 32'hEA752DFE
`define SBOX1_ELEMENT_199 32'h8B021FA1
`define SBOX1_ELEMENT_200 32'hE5A0CC0F
`define SBOX1_ELEMENT_201 32'hB56F74E8
`define SBOX1_ELEMENT_202 32'h18ACF3D6
`define SBOX1_ELEMENT_203 32'hCE89E299
`define SBOX1_ELEMENT_204 32'hB4A84FE0
`define SBOX1_ELEMENT_205 32'hFD13E0B7
`define SBOX1_ELEMENT_206 32'h7CC43B81
`define SBOX1_ELEMENT_207 32'hD2ADA8D9
`define SBOX1_ELEMENT_208 32'h165FA266
`define SBOX1_ELEMENT_209 32'h80957705
`define SBOX1_ELEMENT_210 32'h93CC7314
`define SBOX1_ELEMENT_211 32'h211A1477
`define SBOX1_ELEMENT_212 32'hE6AD2065
`define SBOX1_ELEMENT_213 32'h77B5FA86
`define SBOX1_ELEMENT_214 32'hC75442F5
`define SBOX1_ELEMENT_215 32'hFB9D35CF
`define SBOX1_ELEMENT_216 32'hEBCDAF0C
`define SBOX1_ELEMENT_217 32'h7B3E89A0
`define SBOX1_ELEMENT_218 32'hD6411BD3
`define SBOX1_ELEMENT_219 32'hAE1E7E49
`define SBOX1_ELEMENT_220 32'h00250E2D
`define SBOX1_ELEMENT_221 32'h2071B35E
`define SBOX1_ELEMENT_222 32'h226800BB
`define SBOX1_ELEMENT_223 32'h57B8E0AF
`define SBOX1_ELEMENT_224 32'h2464369B
`define SBOX1_ELEMENT_225 32'hF009B91E
`define SBOX1_ELEMENT_226 32'h5563911D
`define SBOX1_ELEMENT_227 32'h59DFA6AA
`define SBOX1_ELEMENT_228 32'h78C14389
`define SBOX1_ELEMENT_229 32'hD95A537F
`define SBOX1_ELEMENT_230 32'h207D5BA2
`define SBOX1_ELEMENT_231 32'h02E5B9C5
`define SBOX1_ELEMENT_232 32'h83260376
`define SBOX1_ELEMENT_233 32'h6295CFA9
`define SBOX1_ELEMENT_234 32'h11C81968
`define SBOX1_ELEMENT_235 32'h4E734A41
`define SBOX1_ELEMENT_236 32'hB3472DCA
`define SBOX1_ELEMENT_237 32'h7B14A94A
`define SBOX1_ELEMENT_238 32'h1B510052
`define SBOX1_ELEMENT_239 32'h9A532915
`define SBOX1_ELEMENT_240 32'hD60F573F
`define SBOX1_ELEMENT_241 32'hBC9BC6E4
`define SBOX1_ELEMENT_242 32'h2B60A476
`define SBOX1_ELEMENT_243 32'h81E67400
`define SBOX1_ELEMENT_244 32'h08BA6FB5
`define SBOX1_ELEMENT_245 32'h571BE91F
`define SBOX1_ELEMENT_246 32'hF296EC6B
`define SBOX1_ELEMENT_247 32'h2A0DD915
`define SBOX1_ELEMENT_248 32'hB6636521
`define SBOX1_ELEMENT_249 32'hE7B9F9B6
`define SBOX1_ELEMENT_250 32'hFF34052E
`define SBOX1_ELEMENT_251 32'hC5855664
`define SBOX1_ELEMENT_252 32'h53B02D5D
`define SBOX1_ELEMENT_253 32'hA99F8FA1
`define SBOX1_ELEMENT_254 32'h08BA4799
`define SBOX1_ELEMENT_255 32'h6E85076A

//SBox2 Macro's Values
`define SBOX2_ELEMENT_000 32'h4B7A70E9
`define SBOX2_ELEMENT_001 32'hB5B32944
`define SBOX2_ELEMENT_002 32'hDB75092E
`define SBOX2_ELEMENT_003 32'hC4192623
`define SBOX2_ELEMENT_004 32'hAD6EA6B0
`define SBOX2_ELEMENT_005 32'h49A7DF7D
`define SBOX2_ELEMENT_006 32'h9CEE60B8
`define SBOX2_ELEMENT_007 32'h8FEDB266
`define SBOX2_ELEMENT_008 32'hECAA8C71
`define SBOX2_ELEMENT_009 32'h699A17FF
`define SBOX2_ELEMENT_010 32'h5664526C
`define SBOX2_ELEMENT_011 32'hC2B19EE1
`define SBOX2_ELEMENT_012 32'h193602A5
`define SBOX2_ELEMENT_013 32'h75094C29
`define SBOX2_ELEMENT_014 32'hA0591340
`define SBOX2_ELEMENT_015 32'hE4183A3E
`define SBOX2_ELEMENT_016 32'h3F54989A
`define SBOX2_ELEMENT_017 32'h5B429D65
`define SBOX2_ELEMENT_018 32'h6B8FE4D6
`define SBOX2_ELEMENT_019 32'h99F73FD6
`define SBOX2_ELEMENT_020 32'hA1D29C07
`define SBOX2_ELEMENT_021 32'hEFE830F5
`define SBOX2_ELEMENT_022 32'h4D2D38E6
`define SBOX2_ELEMENT_023 32'hF0255DC1
`define SBOX2_ELEMENT_024 32'h4CDD2086
`define SBOX2_ELEMENT_025 32'h8470EB26
`define SBOX2_ELEMENT_026 32'h6382E9C6
`define SBOX2_ELEMENT_027 32'h021ECC5E
`define SBOX2_ELEMENT_028 32'h09686B3F
`define SBOX2_ELEMENT_029 32'h3EBAEFC9
`define SBOX2_ELEMENT_030 32'h3C971814
`define SBOX2_ELEMENT_031 32'h6B6A70A1
`define SBOX2_ELEMENT_032 32'h687F3584
`define SBOX2_ELEMENT_033 32'h52A0E286
`define SBOX2_ELEMENT_034 32'hB79C5305
`define SBOX2_ELEMENT_035 32'hAA500737
`define SBOX2_ELEMENT_036 32'h3E07841C
`define SBOX2_ELEMENT_037 32'h7FDEAE5C
`define SBOX2_ELEMENT_038 32'h8E7D44EC
`define SBOX2_ELEMENT_039 32'h5716F2B8
`define SBOX2_ELEMENT_040 32'hB03ADA37
`define SBOX2_ELEMENT_041 32'hF0500C0D
`define SBOX2_ELEMENT_042 32'hF01C1F04
`define SBOX2_ELEMENT_043 32'h0200B3FF
`define SBOX2_ELEMENT_044 32'hAE0CF51A
`define SBOX2_ELEMENT_045 32'h3CB574B2
`define SBOX2_ELEMENT_046 32'h25837A58
`define SBOX2_ELEMENT_047 32'hDC0921BD
`define SBOX2_ELEMENT_048 32'hD19113F9
`define SBOX2_ELEMENT_049 32'h7CA92FF6
`define SBOX2_ELEMENT_050 32'h94324773
`define SBOX2_ELEMENT_051 32'h22F54701
`define SBOX2_ELEMENT_052 32'h3AE5E581
`define SBOX2_ELEMENT_053 32'h37C2DADC
`define SBOX2_ELEMENT_054 32'hC8B57634
`define SBOX2_ELEMENT_055 32'h9AF3DDA7
`define SBOX2_ELEMENT_056 32'hA9446146
`define SBOX2_ELEMENT_057 32'h0FD0030E
`define SBOX2_ELEMENT_058 32'hECC8C73E
`define SBOX2_ELEMENT_059 32'hA4751E41
`define SBOX2_ELEMENT_060 32'hE238CD99
`define SBOX2_ELEMENT_061 32'h3BEA0E2F
`define SBOX2_ELEMENT_062 32'h3280BBA1
`define SBOX2_ELEMENT_063 32'h183EB331
`define SBOX2_ELEMENT_064 32'h4E548B38
`define SBOX2_ELEMENT_065 32'h4F6DB908
`define SBOX2_ELEMENT_066 32'h6F420D03
`define SBOX2_ELEMENT_067 32'hF60A04BF
`define SBOX2_ELEMENT_068 32'h2CB81290
`define SBOX2_ELEMENT_069 32'h24977C79
`define SBOX2_ELEMENT_070 32'h5679B072
`define SBOX2_ELEMENT_071 32'hBCAF89AF
`define SBOX2_ELEMENT_072 32'hDE9A771F
`define SBOX2_ELEMENT_073 32'hD9930810
`define SBOX2_ELEMENT_074 32'hB38BAE12
`define SBOX2_ELEMENT_075 32'hDCCF3F2E
`define SBOX2_ELEMENT_076 32'h5512721F
`define SBOX2_ELEMENT_077 32'h2E6B7124
`define SBOX2_ELEMENT_078 32'h501ADDE6
`define SBOX2_ELEMENT_079 32'h9F84CD87
`define SBOX2_ELEMENT_080 32'h7A584718
`define SBOX2_ELEMENT_081 32'h7408DA17
`define SBOX2_ELEMENT_082 32'hBC9F9ABC
`define SBOX2_ELEMENT_083 32'hE94B7D8C
`define SBOX2_ELEMENT_084 32'hEC7AEC3A
`define SBOX2_ELEMENT_085 32'hDB851DFA
`define SBOX2_ELEMENT_086 32'h63094366
`define SBOX2_ELEMENT_087 32'hC464C3D2
`define SBOX2_ELEMENT_088 32'hEF1C1847
`define SBOX2_ELEMENT_089 32'h3215D908
`define SBOX2_ELEMENT_090 32'hDD433B37
`define SBOX2_ELEMENT_091 32'h24C2BA16
`define SBOX2_ELEMENT_092 32'h12A14D43
`define SBOX2_ELEMENT_093 32'h2A65C451
`define SBOX2_ELEMENT_094 32'h50940002
`define SBOX2_ELEMENT_095 32'h133AE4DD
`define SBOX2_ELEMENT_096 32'h71DFF89E
`define SBOX2_ELEMENT_097 32'h10314E55
`define SBOX2_ELEMENT_098 32'h81AC77D6
`define SBOX2_ELEMENT_099 32'h5F11199B
`define SBOX2_ELEMENT_100 32'h043556F1
`define SBOX2_ELEMENT_101 32'hD7A3C76B
`define SBOX2_ELEMENT_102 32'h3C11183B
`define SBOX2_ELEMENT_103 32'h5924A509
`define SBOX2_ELEMENT_104 32'hF28FE6ED
`define SBOX2_ELEMENT_105 32'h97F1FBFA
`define SBOX2_ELEMENT_106 32'h9EBABF2C
`define SBOX2_ELEMENT_107 32'h1E153C6E
`define SBOX2_ELEMENT_108 32'h86E34570
`define SBOX2_ELEMENT_109 32'hEAE96FB1
`define SBOX2_ELEMENT_110 32'h860E5E0A
`define SBOX2_ELEMENT_111 32'h5A3E2AB3
`define SBOX2_ELEMENT_112 32'h771FE71C
`define SBOX2_ELEMENT_113 32'h4E3D06FA
`define SBOX2_ELEMENT_114 32'h2965DCB9
`define SBOX2_ELEMENT_115 32'h99E71D0F
`define SBOX2_ELEMENT_116 32'h803E89D6
`define SBOX2_ELEMENT_117 32'h5266C825
`define SBOX2_ELEMENT_118 32'h2E4CC978
`define SBOX2_ELEMENT_119 32'h9C10B36A
`define SBOX2_ELEMENT_120 32'hC6150EBA
`define SBOX2_ELEMENT_121 32'h94E2EA78
`define SBOX2_ELEMENT_122 32'hA5FC3C53
`define SBOX2_ELEMENT_123 32'h1E0A2DF4
`define SBOX2_ELEMENT_124 32'hF2F74EA7
`define SBOX2_ELEMENT_125 32'h361D2B3D
`define SBOX2_ELEMENT_126 32'h1939260F
`define SBOX2_ELEMENT_127 32'h19C27960
`define SBOX2_ELEMENT_128 32'h5223A708
`define SBOX2_ELEMENT_129 32'hF71312B6
`define SBOX2_ELEMENT_130 32'hEBADFE6E
`define SBOX2_ELEMENT_131 32'hEAC31F66
`define SBOX2_ELEMENT_132 32'hE3BC4595
`define SBOX2_ELEMENT_133 32'hA67BC883
`define SBOX2_ELEMENT_134 32'hB17F37D1
`define SBOX2_ELEMENT_135 32'h018CFF28
`define SBOX2_ELEMENT_136 32'hC332DDEF
`define SBOX2_ELEMENT_137 32'hBE6C5AA5
`define SBOX2_ELEMENT_138 32'h65582185
`define SBOX2_ELEMENT_139 32'h68AB9802
`define SBOX2_ELEMENT_140 32'hEECEA50F
`define SBOX2_ELEMENT_141 32'hDB2F953B
`define SBOX2_ELEMENT_142 32'h2AEF7DAD
`define SBOX2_ELEMENT_143 32'h5B6E2F84
`define SBOX2_ELEMENT_144 32'h1521B628
`define SBOX2_ELEMENT_145 32'h29076170
`define SBOX2_ELEMENT_146 32'hECDD4775
`define SBOX2_ELEMENT_147 32'h619F1510
`define SBOX2_ELEMENT_148 32'h13CCA830
`define SBOX2_ELEMENT_149 32'hEB61BD96
`define SBOX2_ELEMENT_150 32'h0334FE1E
`define SBOX2_ELEMENT_151 32'hAA0363CF
`define SBOX2_ELEMENT_152 32'hB5735C90
`define SBOX2_ELEMENT_153 32'h4C70A239
`define SBOX2_ELEMENT_154 32'hD59E9E0B
`define SBOX2_ELEMENT_155 32'hCBAADE14
`define SBOX2_ELEMENT_156 32'hEECC86BC
`define SBOX2_ELEMENT_157 32'h60622CA7
`define SBOX2_ELEMENT_158 32'h9CAB5CAB
`define SBOX2_ELEMENT_159 32'hB2F3846E
`define SBOX2_ELEMENT_160 32'h648B1EAF
`define SBOX2_ELEMENT_161 32'h19BDF0CA
`define SBOX2_ELEMENT_162 32'hA02369B9
`define SBOX2_ELEMENT_163 32'h655ABB50
`define SBOX2_ELEMENT_164 32'h40685A32
`define SBOX2_ELEMENT_165 32'h3C2AB4B3
`define SBOX2_ELEMENT_166 32'h319EE9D5
`define SBOX2_ELEMENT_167 32'hC021B8F7
`define SBOX2_ELEMENT_168 32'h9B540B19
`define SBOX2_ELEMENT_169 32'h875FA099
`define SBOX2_ELEMENT_170 32'h95F7997E
`define SBOX2_ELEMENT_171 32'h623D7DA8
`define SBOX2_ELEMENT_172 32'hF837889A
`define SBOX2_ELEMENT_173 32'h97E32D77
`define SBOX2_ELEMENT_174 32'h11ED935F
`define SBOX2_ELEMENT_175 32'h16681281
`define SBOX2_ELEMENT_176 32'h0E358829
`define SBOX2_ELEMENT_177 32'hC7E61FD6
`define SBOX2_ELEMENT_178 32'h96DEDFA1
`define SBOX2_ELEMENT_179 32'h7858BA99
`define SBOX2_ELEMENT_180 32'h57F584A5
`define SBOX2_ELEMENT_181 32'h1B227263
`define SBOX2_ELEMENT_182 32'h9B83C3FF
`define SBOX2_ELEMENT_183 32'h1AC24696
`define SBOX2_ELEMENT_184 32'hCDB30AEB
`define SBOX2_ELEMENT_185 32'h532E3054
`define SBOX2_ELEMENT_186 32'h8FD948E4
`define SBOX2_ELEMENT_187 32'h6DBC3128
`define SBOX2_ELEMENT_188 32'h58EBF2EF
`define SBOX2_ELEMENT_189 32'h34C6FFEA
`define SBOX2_ELEMENT_190 32'hFE28ED61
`define SBOX2_ELEMENT_191 32'hEE7C3C73
`define SBOX2_ELEMENT_192 32'h5D4A14D9
`define SBOX2_ELEMENT_193 32'hE864B7E3
`define SBOX2_ELEMENT_194 32'h42105D14
`define SBOX2_ELEMENT_195 32'h203E13E0
`define SBOX2_ELEMENT_196 32'h45EEE2B6
`define SBOX2_ELEMENT_197 32'hA3AAABEA
`define SBOX2_ELEMENT_198 32'hDB6C4F15
`define SBOX2_ELEMENT_199 32'hFACB4FD0
`define SBOX2_ELEMENT_200 32'hC742F442
`define SBOX2_ELEMENT_201 32'hEF6ABBB5
`define SBOX2_ELEMENT_202 32'h654F3B1D
`define SBOX2_ELEMENT_203 32'h41CD2105
`define SBOX2_ELEMENT_204 32'hD81E799E
`define SBOX2_ELEMENT_205 32'h86854DC7
`define SBOX2_ELEMENT_206 32'hE44B476A
`define SBOX2_ELEMENT_207 32'h3D816250
`define SBOX2_ELEMENT_208 32'hCF62A1F2
`define SBOX2_ELEMENT_209 32'h5B8D2646
`define SBOX2_ELEMENT_210 32'hFC8883A0
`define SBOX2_ELEMENT_211 32'hC1C7B6A3
`define SBOX2_ELEMENT_212 32'h7F1524C3
`define SBOX2_ELEMENT_213 32'h69CB7492
`define SBOX2_ELEMENT_214 32'h47848A0B
`define SBOX2_ELEMENT_215 32'h5692B285
`define SBOX2_ELEMENT_216 32'h095BBF00
`define SBOX2_ELEMENT_217 32'hAD19489D
`define SBOX2_ELEMENT_218 32'h1462B174
`define SBOX2_ELEMENT_219 32'h23820E00
`define SBOX2_ELEMENT_220 32'h58428D2A
`define SBOX2_ELEMENT_221 32'h0C55F5EA
`define SBOX2_ELEMENT_222 32'h1DADF43E
`define SBOX2_ELEMENT_223 32'h233F7061
`define SBOX2_ELEMENT_224 32'h3372F092
`define SBOX2_ELEMENT_225 32'h8D937E41
`define SBOX2_ELEMENT_226 32'hD65FECF1
`define SBOX2_ELEMENT_227 32'h6C223BDB
`define SBOX2_ELEMENT_228 32'h7CDE3759
`define SBOX2_ELEMENT_229 32'hCBEE7460
`define SBOX2_ELEMENT_230 32'h4085F2A7
`define SBOX2_ELEMENT_231 32'hCE77326E
`define SBOX2_ELEMENT_232 32'hA6078084
`define SBOX2_ELEMENT_233 32'h19F8509E
`define SBOX2_ELEMENT_234 32'hE8EFD855
`define SBOX2_ELEMENT_235 32'h61D99735
`define SBOX2_ELEMENT_236 32'hA969A7AA
`define SBOX2_ELEMENT_237 32'hC50C06C2
`define SBOX2_ELEMENT_238 32'h5A04ABFC
`define SBOX2_ELEMENT_239 32'h800BCADC
`define SBOX2_ELEMENT_240 32'h9E447A2E
`define SBOX2_ELEMENT_241 32'hC3453484
`define SBOX2_ELEMENT_242 32'hFDD56705
`define SBOX2_ELEMENT_243 32'h0E1E9EC9
`define SBOX2_ELEMENT_244 32'hDB73DBD3
`define SBOX2_ELEMENT_245 32'h105588CD
`define SBOX2_ELEMENT_246 32'h675FDA79
`define SBOX2_ELEMENT_247 32'hE3674340
`define SBOX2_ELEMENT_248 32'hC5C43465
`define SBOX2_ELEMENT_249 32'h713E38D8
`define SBOX2_ELEMENT_250 32'h3D28F89E
`define SBOX2_ELEMENT_251 32'hF16DFF20
`define SBOX2_ELEMENT_252 32'h153E21E7
`define SBOX2_ELEMENT_253 32'h8FB03D4A
`define SBOX2_ELEMENT_254 32'hE6E39F2B
`define SBOX2_ELEMENT_255 32'hDB83ADF7
