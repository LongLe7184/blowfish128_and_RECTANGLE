//-----------------------------------------------------------
// Function: Blowfish-128's S-Boxes
//-----------------------------------------------------------
// Author	: Long Le, Manh Nguyen
// Date  	: Feb-5th, 2025
// Description	: Contains 2 Substitution Boxes, each has 256 elements 32-bit
//-----------------------------------------------------------

`include "blowfish128_DEF.vh"

//Include Guards - avoid declare multiple times
`ifndef BLOWFISH128_SBOX
`define BLOWFISH128_SBOX

module blowfish128_sbox1(
	input [7:0] sbox_in,
	output reg [31:0] sbox_out
	);

	always @(*) begin
		case (sbox_in[7:0])
			8'h00: sbox_out = `SBOX1_ELEMENT_000;
			8'h01: sbox_out = `SBOX1_ELEMENT_001;
			8'h02: sbox_out = `SBOX1_ELEMENT_002;
			8'h03: sbox_out = `SBOX1_ELEMENT_003;
			8'h04: sbox_out = `SBOX1_ELEMENT_004;
			8'h05: sbox_out = `SBOX1_ELEMENT_005;
			8'h06: sbox_out = `SBOX1_ELEMENT_006;
			8'h07: sbox_out = `SBOX1_ELEMENT_007;
			8'h08: sbox_out = `SBOX1_ELEMENT_008;
			8'h09: sbox_out = `SBOX1_ELEMENT_009;
			8'h0A: sbox_out = `SBOX1_ELEMENT_010;
			8'h0B: sbox_out = `SBOX1_ELEMENT_011;
			8'h0C: sbox_out = `SBOX1_ELEMENT_012;
			8'h0D: sbox_out = `SBOX1_ELEMENT_013;
			8'h0E: sbox_out = `SBOX1_ELEMENT_014;
			8'h0F: sbox_out = `SBOX1_ELEMENT_015;
			8'h10: sbox_out = `SBOX1_ELEMENT_016;
			8'h11: sbox_out = `SBOX1_ELEMENT_017;
			8'h12: sbox_out = `SBOX1_ELEMENT_018;
			8'h13: sbox_out = `SBOX1_ELEMENT_019;
			8'h14: sbox_out = `SBOX1_ELEMENT_020;
			8'h15: sbox_out = `SBOX1_ELEMENT_021;
			8'h16: sbox_out = `SBOX1_ELEMENT_022;
			8'h17: sbox_out = `SBOX1_ELEMENT_023;
			8'h18: sbox_out = `SBOX1_ELEMENT_024;
			8'h19: sbox_out = `SBOX1_ELEMENT_025;
			8'h1A: sbox_out = `SBOX1_ELEMENT_026;
			8'h1B: sbox_out = `SBOX1_ELEMENT_027;
			8'h1C: sbox_out = `SBOX1_ELEMENT_028;
			8'h1D: sbox_out = `SBOX1_ELEMENT_029;
			8'h1E: sbox_out = `SBOX1_ELEMENT_030;
			8'h1F: sbox_out = `SBOX1_ELEMENT_031;
			8'h20: sbox_out = `SBOX1_ELEMENT_032;
			8'h21: sbox_out = `SBOX1_ELEMENT_033;
			8'h22: sbox_out = `SBOX1_ELEMENT_034;
			8'h23: sbox_out = `SBOX1_ELEMENT_035;
			8'h24: sbox_out = `SBOX1_ELEMENT_036;
			8'h25: sbox_out = `SBOX1_ELEMENT_037;
			8'h26: sbox_out = `SBOX1_ELEMENT_038;
			8'h27: sbox_out = `SBOX1_ELEMENT_039;
			8'h28: sbox_out = `SBOX1_ELEMENT_040;
			8'h29: sbox_out = `SBOX1_ELEMENT_041;
			8'h2A: sbox_out = `SBOX1_ELEMENT_042;
			8'h2B: sbox_out = `SBOX1_ELEMENT_043;
			8'h2C: sbox_out = `SBOX1_ELEMENT_044;
			8'h2D: sbox_out = `SBOX1_ELEMENT_045;
			8'h2E: sbox_out = `SBOX1_ELEMENT_046;
			8'h2F: sbox_out = `SBOX1_ELEMENT_047;
			8'h30: sbox_out = `SBOX1_ELEMENT_048;
			8'h31: sbox_out = `SBOX1_ELEMENT_049;
			8'h32: sbox_out = `SBOX1_ELEMENT_050;
			8'h33: sbox_out = `SBOX1_ELEMENT_051;
			8'h34: sbox_out = `SBOX1_ELEMENT_052;
			8'h35: sbox_out = `SBOX1_ELEMENT_053;
			8'h36: sbox_out = `SBOX1_ELEMENT_054;
			8'h37: sbox_out = `SBOX1_ELEMENT_055;
			8'h38: sbox_out = `SBOX1_ELEMENT_056;
			8'h39: sbox_out = `SBOX1_ELEMENT_057;
			8'h3A: sbox_out = `SBOX1_ELEMENT_058;
			8'h3B: sbox_out = `SBOX1_ELEMENT_059;
			8'h3C: sbox_out = `SBOX1_ELEMENT_060;
			8'h3D: sbox_out = `SBOX1_ELEMENT_061;
			8'h3E: sbox_out = `SBOX1_ELEMENT_062;
			8'h3F: sbox_out = `SBOX1_ELEMENT_063;
			8'h40: sbox_out = `SBOX1_ELEMENT_064;
			8'h41: sbox_out = `SBOX1_ELEMENT_065;
			8'h42: sbox_out = `SBOX1_ELEMENT_066;
			8'h43: sbox_out = `SBOX1_ELEMENT_067;
			8'h44: sbox_out = `SBOX1_ELEMENT_068;
			8'h45: sbox_out = `SBOX1_ELEMENT_069;
			8'h46: sbox_out = `SBOX1_ELEMENT_070;
			8'h47: sbox_out = `SBOX1_ELEMENT_071;
			8'h48: sbox_out = `SBOX1_ELEMENT_072;
			8'h49: sbox_out = `SBOX1_ELEMENT_073;
			8'h4A: sbox_out = `SBOX1_ELEMENT_074;
			8'h4B: sbox_out = `SBOX1_ELEMENT_075;
			8'h4C: sbox_out = `SBOX1_ELEMENT_076;
			8'h4D: sbox_out = `SBOX1_ELEMENT_077;
			8'h4E: sbox_out = `SBOX1_ELEMENT_078;
			8'h4F: sbox_out = `SBOX1_ELEMENT_079;
			8'h50: sbox_out = `SBOX1_ELEMENT_080;
			8'h51: sbox_out = `SBOX1_ELEMENT_081;
			8'h52: sbox_out = `SBOX1_ELEMENT_082;
			8'h53: sbox_out = `SBOX1_ELEMENT_083;
			8'h54: sbox_out = `SBOX1_ELEMENT_084;
			8'h55: sbox_out = `SBOX1_ELEMENT_085;
			8'h56: sbox_out = `SBOX1_ELEMENT_086;
			8'h57: sbox_out = `SBOX1_ELEMENT_087;
			8'h58: sbox_out = `SBOX1_ELEMENT_088;
			8'h59: sbox_out = `SBOX1_ELEMENT_089;
			8'h5A: sbox_out = `SBOX1_ELEMENT_090;
			8'h5B: sbox_out = `SBOX1_ELEMENT_091;
			8'h5C: sbox_out = `SBOX1_ELEMENT_092;
			8'h5D: sbox_out = `SBOX1_ELEMENT_093;
			8'h5E: sbox_out = `SBOX1_ELEMENT_094;
			8'h5F: sbox_out = `SBOX1_ELEMENT_095;
			8'h60: sbox_out = `SBOX1_ELEMENT_096;
			8'h61: sbox_out = `SBOX1_ELEMENT_097;
			8'h62: sbox_out = `SBOX1_ELEMENT_098;
			8'h63: sbox_out = `SBOX1_ELEMENT_099;
			8'h64: sbox_out = `SBOX1_ELEMENT_100;
			8'h65: sbox_out = `SBOX1_ELEMENT_101;
			8'h66: sbox_out = `SBOX1_ELEMENT_102;
			8'h67: sbox_out = `SBOX1_ELEMENT_103;
			8'h68: sbox_out = `SBOX1_ELEMENT_104;
			8'h69: sbox_out = `SBOX1_ELEMENT_105;
			8'h6A: sbox_out = `SBOX1_ELEMENT_106;
			8'h6B: sbox_out = `SBOX1_ELEMENT_107;
			8'h6C: sbox_out = `SBOX1_ELEMENT_108;
			8'h6D: sbox_out = `SBOX1_ELEMENT_109;
			8'h6E: sbox_out = `SBOX1_ELEMENT_110;
			8'h6F: sbox_out = `SBOX1_ELEMENT_111;
			8'h70: sbox_out = `SBOX1_ELEMENT_112;
			8'h71: sbox_out = `SBOX1_ELEMENT_113;
			8'h72: sbox_out = `SBOX1_ELEMENT_114;
			8'h73: sbox_out = `SBOX1_ELEMENT_115;
			8'h74: sbox_out = `SBOX1_ELEMENT_116;
			8'h75: sbox_out = `SBOX1_ELEMENT_117;
			8'h76: sbox_out = `SBOX1_ELEMENT_118;
			8'h77: sbox_out = `SBOX1_ELEMENT_119;
			8'h78: sbox_out = `SBOX1_ELEMENT_120;
			8'h79: sbox_out = `SBOX1_ELEMENT_121;
			8'h7A: sbox_out = `SBOX1_ELEMENT_122;
			8'h7B: sbox_out = `SBOX1_ELEMENT_123;
			8'h7C: sbox_out = `SBOX1_ELEMENT_124;
			8'h7D: sbox_out = `SBOX1_ELEMENT_125;
			8'h7E: sbox_out = `SBOX1_ELEMENT_126;
			8'h7F: sbox_out = `SBOX1_ELEMENT_127;
			8'h80: sbox_out = `SBOX1_ELEMENT_128;
			8'h81: sbox_out = `SBOX1_ELEMENT_129;
			8'h82: sbox_out = `SBOX1_ELEMENT_130;
			8'h83: sbox_out = `SBOX1_ELEMENT_131;
			8'h84: sbox_out = `SBOX1_ELEMENT_132;
			8'h85: sbox_out = `SBOX1_ELEMENT_133;
			8'h86: sbox_out = `SBOX1_ELEMENT_134;
			8'h87: sbox_out = `SBOX1_ELEMENT_135;
			8'h88: sbox_out = `SBOX1_ELEMENT_136;
			8'h89: sbox_out = `SBOX1_ELEMENT_137;
			8'h8A: sbox_out = `SBOX1_ELEMENT_138;
			8'h8B: sbox_out = `SBOX1_ELEMENT_139;
			8'h8C: sbox_out = `SBOX1_ELEMENT_140;
			8'h8D: sbox_out = `SBOX1_ELEMENT_141;
			8'h8E: sbox_out = `SBOX1_ELEMENT_142;
			8'h8F: sbox_out = `SBOX1_ELEMENT_143;
			8'h90: sbox_out = `SBOX1_ELEMENT_144;
			8'h91: sbox_out = `SBOX1_ELEMENT_145;
			8'h92: sbox_out = `SBOX1_ELEMENT_146;
			8'h93: sbox_out = `SBOX1_ELEMENT_147;
			8'h94: sbox_out = `SBOX1_ELEMENT_148;
			8'h95: sbox_out = `SBOX1_ELEMENT_149;
			8'h96: sbox_out = `SBOX1_ELEMENT_150;
			8'h97: sbox_out = `SBOX1_ELEMENT_151;
			8'h98: sbox_out = `SBOX1_ELEMENT_152;
			8'h99: sbox_out = `SBOX1_ELEMENT_153;
			8'h9A: sbox_out = `SBOX1_ELEMENT_154;
			8'h9B: sbox_out = `SBOX1_ELEMENT_155;
			8'h9C: sbox_out = `SBOX1_ELEMENT_156;
			8'h9D: sbox_out = `SBOX1_ELEMENT_157;
			8'h9E: sbox_out = `SBOX1_ELEMENT_158;
			8'h9F: sbox_out = `SBOX1_ELEMENT_159;
			8'hA0: sbox_out = `SBOX1_ELEMENT_160;
			8'hA1: sbox_out = `SBOX1_ELEMENT_161;
			8'hA2: sbox_out = `SBOX1_ELEMENT_162;
			8'hA3: sbox_out = `SBOX1_ELEMENT_163;
			8'hA4: sbox_out = `SBOX1_ELEMENT_164;
			8'hA5: sbox_out = `SBOX1_ELEMENT_165;
			8'hA6: sbox_out = `SBOX1_ELEMENT_166;
			8'hA7: sbox_out = `SBOX1_ELEMENT_167;
			8'hA8: sbox_out = `SBOX1_ELEMENT_168;
			8'hA9: sbox_out = `SBOX1_ELEMENT_169;
			8'hAA: sbox_out = `SBOX1_ELEMENT_170;
			8'hAB: sbox_out = `SBOX1_ELEMENT_171;
			8'hAC: sbox_out = `SBOX1_ELEMENT_172;
			8'hAD: sbox_out = `SBOX1_ELEMENT_173;
			8'hAE: sbox_out = `SBOX1_ELEMENT_174;
			8'hAF: sbox_out = `SBOX1_ELEMENT_175;
			8'hB0: sbox_out = `SBOX1_ELEMENT_176;
			8'hB1: sbox_out = `SBOX1_ELEMENT_177;
			8'hB2: sbox_out = `SBOX1_ELEMENT_178;
			8'hB3: sbox_out = `SBOX1_ELEMENT_179;
			8'hB4: sbox_out = `SBOX1_ELEMENT_180;
			8'hB5: sbox_out = `SBOX1_ELEMENT_181;
			8'hB6: sbox_out = `SBOX1_ELEMENT_182;
			8'hB7: sbox_out = `SBOX1_ELEMENT_183;
			8'hB8: sbox_out = `SBOX1_ELEMENT_184;
			8'hB9: sbox_out = `SBOX1_ELEMENT_185;
			8'hBA: sbox_out = `SBOX1_ELEMENT_186;
			8'hBB: sbox_out = `SBOX1_ELEMENT_187;
			8'hBC: sbox_out = `SBOX1_ELEMENT_188;
			8'hBD: sbox_out = `SBOX1_ELEMENT_189;
			8'hBE: sbox_out = `SBOX1_ELEMENT_190;
			8'hBF: sbox_out = `SBOX1_ELEMENT_191;
			8'hC0: sbox_out = `SBOX1_ELEMENT_192;
			8'hC1: sbox_out = `SBOX1_ELEMENT_193;
			8'hC2: sbox_out = `SBOX1_ELEMENT_194;
			8'hC3: sbox_out = `SBOX1_ELEMENT_195;
			8'hC4: sbox_out = `SBOX1_ELEMENT_196;
			8'hC5: sbox_out = `SBOX1_ELEMENT_197;
			8'hC6: sbox_out = `SBOX1_ELEMENT_198;
			8'hC7: sbox_out = `SBOX1_ELEMENT_199;
			8'hC8: sbox_out = `SBOX1_ELEMENT_200;
			8'hC9: sbox_out = `SBOX1_ELEMENT_201;
			8'hCA: sbox_out = `SBOX1_ELEMENT_202;
			8'hCB: sbox_out = `SBOX1_ELEMENT_203;
			8'hCC: sbox_out = `SBOX1_ELEMENT_204;
			8'hCD: sbox_out = `SBOX1_ELEMENT_205;
			8'hCE: sbox_out = `SBOX1_ELEMENT_206;
			8'hCF: sbox_out = `SBOX1_ELEMENT_207;
			8'hD0: sbox_out = `SBOX1_ELEMENT_208;
			8'hD1: sbox_out = `SBOX1_ELEMENT_209;
			8'hD2: sbox_out = `SBOX1_ELEMENT_210;
			8'hD3: sbox_out = `SBOX1_ELEMENT_211;
			8'hD4: sbox_out = `SBOX1_ELEMENT_212;
			8'hD5: sbox_out = `SBOX1_ELEMENT_213;
			8'hD6: sbox_out = `SBOX1_ELEMENT_214;
			8'hD7: sbox_out = `SBOX1_ELEMENT_215;
			8'hD8: sbox_out = `SBOX1_ELEMENT_216;
			8'hD9: sbox_out = `SBOX1_ELEMENT_217;
			8'hDA: sbox_out = `SBOX1_ELEMENT_218;
			8'hDB: sbox_out = `SBOX1_ELEMENT_219;
			8'hDC: sbox_out = `SBOX1_ELEMENT_220;
			8'hDD: sbox_out = `SBOX1_ELEMENT_221;
			8'hDE: sbox_out = `SBOX1_ELEMENT_222;
			8'hDF: sbox_out = `SBOX1_ELEMENT_223;
			8'hE0: sbox_out = `SBOX1_ELEMENT_224;
			8'hE1: sbox_out = `SBOX1_ELEMENT_225;
			8'hE2: sbox_out = `SBOX1_ELEMENT_226;
			8'hE3: sbox_out = `SBOX1_ELEMENT_227;
			8'hE4: sbox_out = `SBOX1_ELEMENT_228;
			8'hE5: sbox_out = `SBOX1_ELEMENT_229;
			8'hE6: sbox_out = `SBOX1_ELEMENT_230;
			8'hE7: sbox_out = `SBOX1_ELEMENT_231;
			8'hE8: sbox_out = `SBOX1_ELEMENT_232;
			8'hE9: sbox_out = `SBOX1_ELEMENT_233;
			8'hEA: sbox_out = `SBOX1_ELEMENT_234;
			8'hEB: sbox_out = `SBOX1_ELEMENT_235;
			8'hEC: sbox_out = `SBOX1_ELEMENT_236;
			8'hED: sbox_out = `SBOX1_ELEMENT_237;
			8'hEE: sbox_out = `SBOX1_ELEMENT_238;
			8'hEF: sbox_out = `SBOX1_ELEMENT_239;
			8'hF0: sbox_out = `SBOX1_ELEMENT_240;
			8'hF1: sbox_out = `SBOX1_ELEMENT_241;
			8'hF2: sbox_out = `SBOX1_ELEMENT_242;
			8'hF3: sbox_out = `SBOX1_ELEMENT_243;
			8'hF4: sbox_out = `SBOX1_ELEMENT_244;
			8'hF5: sbox_out = `SBOX1_ELEMENT_245;
			8'hF6: sbox_out = `SBOX1_ELEMENT_246;
			8'hF7: sbox_out = `SBOX1_ELEMENT_247;
			8'hF8: sbox_out = `SBOX1_ELEMENT_248;
			8'hF9: sbox_out = `SBOX1_ELEMENT_249;
			8'hFA: sbox_out = `SBOX1_ELEMENT_250;
			8'hFB: sbox_out = `SBOX1_ELEMENT_251;
			8'hFC: sbox_out = `SBOX1_ELEMENT_252;
			8'hFD: sbox_out = `SBOX1_ELEMENT_253;
			8'hFE: sbox_out = `SBOX1_ELEMENT_254;
			8'hFF: sbox_out = `SBOX1_ELEMENT_255;
			default: sbox_out = 32'h0;
		endcase
	end
endmodule

module blowfish128_sbox2(
	input [7:0] sbox_in,
	output reg [31:0] sbox_out
	);

	always @(*) begin
		case(sbox_in[7:0])
			8'h00: sbox_out = `SBOX2_ELEMENT_000;
			8'h01: sbox_out = `SBOX2_ELEMENT_001;
			8'h02: sbox_out = `SBOX2_ELEMENT_002;
			8'h03: sbox_out = `SBOX2_ELEMENT_003;
			8'h04: sbox_out = `SBOX2_ELEMENT_004;
			8'h05: sbox_out = `SBOX2_ELEMENT_005;
			8'h06: sbox_out = `SBOX2_ELEMENT_006;
			8'h07: sbox_out = `SBOX2_ELEMENT_007;
			8'h08: sbox_out = `SBOX2_ELEMENT_008;
			8'h09: sbox_out = `SBOX2_ELEMENT_009;
			8'h0A: sbox_out = `SBOX2_ELEMENT_010;
			8'h0B: sbox_out = `SBOX2_ELEMENT_011;
			8'h0C: sbox_out = `SBOX2_ELEMENT_012;
			8'h0D: sbox_out = `SBOX2_ELEMENT_013;
			8'h0E: sbox_out = `SBOX2_ELEMENT_014;
			8'h0F: sbox_out = `SBOX2_ELEMENT_015;
			8'h10: sbox_out = `SBOX2_ELEMENT_016;
			8'h11: sbox_out = `SBOX2_ELEMENT_017;
			8'h12: sbox_out = `SBOX2_ELEMENT_018;
			8'h13: sbox_out = `SBOX2_ELEMENT_019;
			8'h14: sbox_out = `SBOX2_ELEMENT_020;
			8'h15: sbox_out = `SBOX2_ELEMENT_021;
			8'h16: sbox_out = `SBOX2_ELEMENT_022;
			8'h17: sbox_out = `SBOX2_ELEMENT_023;
			8'h18: sbox_out = `SBOX2_ELEMENT_024;
			8'h19: sbox_out = `SBOX2_ELEMENT_025;
			8'h1A: sbox_out = `SBOX2_ELEMENT_026;
			8'h1B: sbox_out = `SBOX2_ELEMENT_027;
			8'h1C: sbox_out = `SBOX2_ELEMENT_028;
			8'h1D: sbox_out = `SBOX2_ELEMENT_029;
			8'h1E: sbox_out = `SBOX2_ELEMENT_030;
			8'h1F: sbox_out = `SBOX2_ELEMENT_031;
			8'h20: sbox_out = `SBOX2_ELEMENT_032;
			8'h21: sbox_out = `SBOX2_ELEMENT_033;
			8'h22: sbox_out = `SBOX2_ELEMENT_034;
			8'h23: sbox_out = `SBOX2_ELEMENT_035;
			8'h24: sbox_out = `SBOX2_ELEMENT_036;
			8'h25: sbox_out = `SBOX2_ELEMENT_037;
			8'h26: sbox_out = `SBOX2_ELEMENT_038;
			8'h27: sbox_out = `SBOX2_ELEMENT_039;
			8'h28: sbox_out = `SBOX2_ELEMENT_040;
			8'h29: sbox_out = `SBOX2_ELEMENT_041;
			8'h2A: sbox_out = `SBOX2_ELEMENT_042;
			8'h2B: sbox_out = `SBOX2_ELEMENT_043;
			8'h2C: sbox_out = `SBOX2_ELEMENT_044;
			8'h2D: sbox_out = `SBOX2_ELEMENT_045;
			8'h2E: sbox_out = `SBOX2_ELEMENT_046;
			8'h2F: sbox_out = `SBOX2_ELEMENT_047;
			8'h30: sbox_out = `SBOX2_ELEMENT_048;
			8'h31: sbox_out = `SBOX2_ELEMENT_049;
			8'h32: sbox_out = `SBOX2_ELEMENT_050;
			8'h33: sbox_out = `SBOX2_ELEMENT_051;
			8'h34: sbox_out = `SBOX2_ELEMENT_052;
			8'h35: sbox_out = `SBOX2_ELEMENT_053;
			8'h36: sbox_out = `SBOX2_ELEMENT_054;
			8'h37: sbox_out = `SBOX2_ELEMENT_055;
			8'h38: sbox_out = `SBOX2_ELEMENT_056;
			8'h39: sbox_out = `SBOX2_ELEMENT_057;
			8'h3A: sbox_out = `SBOX2_ELEMENT_058;
			8'h3B: sbox_out = `SBOX2_ELEMENT_059;
			8'h3C: sbox_out = `SBOX2_ELEMENT_060;
			8'h3D: sbox_out = `SBOX2_ELEMENT_061;
			8'h3E: sbox_out = `SBOX2_ELEMENT_062;
			8'h3F: sbox_out = `SBOX2_ELEMENT_063;
			8'h40: sbox_out = `SBOX2_ELEMENT_064;
			8'h41: sbox_out = `SBOX2_ELEMENT_065;
			8'h42: sbox_out = `SBOX2_ELEMENT_066;
			8'h43: sbox_out = `SBOX2_ELEMENT_067;
			8'h44: sbox_out = `SBOX2_ELEMENT_068;
			8'h45: sbox_out = `SBOX2_ELEMENT_069;
			8'h46: sbox_out = `SBOX2_ELEMENT_070;
			8'h47: sbox_out = `SBOX2_ELEMENT_071;
			8'h48: sbox_out = `SBOX2_ELEMENT_072;
			8'h49: sbox_out = `SBOX2_ELEMENT_073;
			8'h4A: sbox_out = `SBOX2_ELEMENT_074;
			8'h4B: sbox_out = `SBOX2_ELEMENT_075;
			8'h4C: sbox_out = `SBOX2_ELEMENT_076;
			8'h4D: sbox_out = `SBOX2_ELEMENT_077;
			8'h4E: sbox_out = `SBOX2_ELEMENT_078;
			8'h4F: sbox_out = `SBOX2_ELEMENT_079;
			8'h50: sbox_out = `SBOX2_ELEMENT_080;
			8'h51: sbox_out = `SBOX2_ELEMENT_081;
			8'h52: sbox_out = `SBOX2_ELEMENT_082;
			8'h53: sbox_out = `SBOX2_ELEMENT_083;
			8'h54: sbox_out = `SBOX2_ELEMENT_084;
			8'h55: sbox_out = `SBOX2_ELEMENT_085;
			8'h56: sbox_out = `SBOX2_ELEMENT_086;
			8'h57: sbox_out = `SBOX2_ELEMENT_087;
			8'h58: sbox_out = `SBOX2_ELEMENT_088;
			8'h59: sbox_out = `SBOX2_ELEMENT_089;
			8'h5A: sbox_out = `SBOX2_ELEMENT_090;
			8'h5B: sbox_out = `SBOX2_ELEMENT_091;
			8'h5C: sbox_out = `SBOX2_ELEMENT_092;
			8'h5D: sbox_out = `SBOX2_ELEMENT_093;
			8'h5E: sbox_out = `SBOX2_ELEMENT_094;
			8'h5F: sbox_out = `SBOX2_ELEMENT_095;
			8'h60: sbox_out = `SBOX2_ELEMENT_096;
			8'h61: sbox_out = `SBOX2_ELEMENT_097;
			8'h62: sbox_out = `SBOX2_ELEMENT_098;
			8'h63: sbox_out = `SBOX2_ELEMENT_099;
			8'h64: sbox_out = `SBOX2_ELEMENT_100;
			8'h65: sbox_out = `SBOX2_ELEMENT_101;
			8'h66: sbox_out = `SBOX2_ELEMENT_102;
			8'h67: sbox_out = `SBOX2_ELEMENT_103;
			8'h68: sbox_out = `SBOX2_ELEMENT_104;
			8'h69: sbox_out = `SBOX2_ELEMENT_105;
			8'h6A: sbox_out = `SBOX2_ELEMENT_106;
			8'h6B: sbox_out = `SBOX2_ELEMENT_107;
			8'h6C: sbox_out = `SBOX2_ELEMENT_108;
			8'h6D: sbox_out = `SBOX2_ELEMENT_109;
			8'h6E: sbox_out = `SBOX2_ELEMENT_110;
			8'h6F: sbox_out = `SBOX2_ELEMENT_111;
			8'h70: sbox_out = `SBOX2_ELEMENT_112;
			8'h71: sbox_out = `SBOX2_ELEMENT_113;
			8'h72: sbox_out = `SBOX2_ELEMENT_114;
			8'h73: sbox_out = `SBOX2_ELEMENT_115;
			8'h74: sbox_out = `SBOX2_ELEMENT_116;
			8'h75: sbox_out = `SBOX2_ELEMENT_117;
			8'h76: sbox_out = `SBOX2_ELEMENT_118;
			8'h77: sbox_out = `SBOX2_ELEMENT_119;
			8'h78: sbox_out = `SBOX2_ELEMENT_120;
			8'h79: sbox_out = `SBOX2_ELEMENT_121;
			8'h7A: sbox_out = `SBOX2_ELEMENT_122;
			8'h7B: sbox_out = `SBOX2_ELEMENT_123;
			8'h7C: sbox_out = `SBOX2_ELEMENT_124;
			8'h7D: sbox_out = `SBOX2_ELEMENT_125;
			8'h7E: sbox_out = `SBOX2_ELEMENT_126;
			8'h7F: sbox_out = `SBOX2_ELEMENT_127;
			8'h80: sbox_out = `SBOX2_ELEMENT_128;
			8'h81: sbox_out = `SBOX2_ELEMENT_129;
			8'h82: sbox_out = `SBOX2_ELEMENT_130;
			8'h83: sbox_out = `SBOX2_ELEMENT_131;
			8'h84: sbox_out = `SBOX2_ELEMENT_132;
			8'h85: sbox_out = `SBOX2_ELEMENT_133;
			8'h86: sbox_out = `SBOX2_ELEMENT_134;
			8'h87: sbox_out = `SBOX2_ELEMENT_135;
			8'h88: sbox_out = `SBOX2_ELEMENT_136;
			8'h89: sbox_out = `SBOX2_ELEMENT_137;
			8'h8A: sbox_out = `SBOX2_ELEMENT_138;
			8'h8B: sbox_out = `SBOX2_ELEMENT_139;
			8'h8C: sbox_out = `SBOX2_ELEMENT_140;
			8'h8D: sbox_out = `SBOX2_ELEMENT_141;
			8'h8E: sbox_out = `SBOX2_ELEMENT_142;
			8'h8F: sbox_out = `SBOX2_ELEMENT_143;
			8'h90: sbox_out = `SBOX2_ELEMENT_144;
			8'h91: sbox_out = `SBOX2_ELEMENT_145;
			8'h92: sbox_out = `SBOX2_ELEMENT_146;
			8'h93: sbox_out = `SBOX2_ELEMENT_147;
			8'h94: sbox_out = `SBOX2_ELEMENT_148;
			8'h95: sbox_out = `SBOX2_ELEMENT_149;
			8'h96: sbox_out = `SBOX2_ELEMENT_150;
			8'h97: sbox_out = `SBOX2_ELEMENT_151;
			8'h98: sbox_out = `SBOX2_ELEMENT_152;
			8'h99: sbox_out = `SBOX2_ELEMENT_153;
			8'h9A: sbox_out = `SBOX2_ELEMENT_154;
			8'h9B: sbox_out = `SBOX2_ELEMENT_155;
			8'h9C: sbox_out = `SBOX2_ELEMENT_156;
			8'h9D: sbox_out = `SBOX2_ELEMENT_157;
			8'h9E: sbox_out = `SBOX2_ELEMENT_158;
			8'h9F: sbox_out = `SBOX2_ELEMENT_159;
			8'hA0: sbox_out = `SBOX2_ELEMENT_160;
			8'hA1: sbox_out = `SBOX2_ELEMENT_161;
			8'hA2: sbox_out = `SBOX2_ELEMENT_162;
			8'hA3: sbox_out = `SBOX2_ELEMENT_163;
			8'hA4: sbox_out = `SBOX2_ELEMENT_164;
			8'hA5: sbox_out = `SBOX2_ELEMENT_165;
			8'hA6: sbox_out = `SBOX2_ELEMENT_166;
			8'hA7: sbox_out = `SBOX2_ELEMENT_167;
			8'hA8: sbox_out = `SBOX2_ELEMENT_168;
			8'hA9: sbox_out = `SBOX2_ELEMENT_169;
			8'hAA: sbox_out = `SBOX2_ELEMENT_170;
			8'hAB: sbox_out = `SBOX2_ELEMENT_171;
			8'hAC: sbox_out = `SBOX2_ELEMENT_172;
			8'hAD: sbox_out = `SBOX2_ELEMENT_173;
			8'hAE: sbox_out = `SBOX2_ELEMENT_174;
			8'hAF: sbox_out = `SBOX2_ELEMENT_175;
			8'hB0: sbox_out = `SBOX2_ELEMENT_176;
			8'hB1: sbox_out = `SBOX2_ELEMENT_177;
			8'hB2: sbox_out = `SBOX2_ELEMENT_178;
			8'hB3: sbox_out = `SBOX2_ELEMENT_179;
			8'hB4: sbox_out = `SBOX2_ELEMENT_180;
			8'hB5: sbox_out = `SBOX2_ELEMENT_181;
			8'hB6: sbox_out = `SBOX2_ELEMENT_182;
			8'hB7: sbox_out = `SBOX2_ELEMENT_183;
			8'hB8: sbox_out = `SBOX2_ELEMENT_184;
			8'hB9: sbox_out = `SBOX2_ELEMENT_185;
			8'hBA: sbox_out = `SBOX2_ELEMENT_186;
			8'hBB: sbox_out = `SBOX2_ELEMENT_187;
			8'hBC: sbox_out = `SBOX2_ELEMENT_188;
			8'hBD: sbox_out = `SBOX2_ELEMENT_189;
			8'hBE: sbox_out = `SBOX2_ELEMENT_190;
			8'hBF: sbox_out = `SBOX2_ELEMENT_191;
			8'hC0: sbox_out = `SBOX2_ELEMENT_192;
			8'hC1: sbox_out = `SBOX2_ELEMENT_193;
			8'hC2: sbox_out = `SBOX2_ELEMENT_194;
			8'hC3: sbox_out = `SBOX2_ELEMENT_195;
			8'hC4: sbox_out = `SBOX2_ELEMENT_196;
			8'hC5: sbox_out = `SBOX2_ELEMENT_197;
			8'hC6: sbox_out = `SBOX2_ELEMENT_198;
			8'hC7: sbox_out = `SBOX2_ELEMENT_199;
			8'hC8: sbox_out = `SBOX2_ELEMENT_200;
			8'hC9: sbox_out = `SBOX2_ELEMENT_201;
			8'hCA: sbox_out = `SBOX2_ELEMENT_202;
			8'hCB: sbox_out = `SBOX2_ELEMENT_203;
			8'hCC: sbox_out = `SBOX2_ELEMENT_204;
			8'hCD: sbox_out = `SBOX2_ELEMENT_205;
			8'hCE: sbox_out = `SBOX2_ELEMENT_206;
			8'hCF: sbox_out = `SBOX2_ELEMENT_207;
			8'hD0: sbox_out = `SBOX2_ELEMENT_208;
			8'hD1: sbox_out = `SBOX2_ELEMENT_209;
			8'hD2: sbox_out = `SBOX2_ELEMENT_210;
			8'hD3: sbox_out = `SBOX2_ELEMENT_211;
			8'hD4: sbox_out = `SBOX2_ELEMENT_212;
			8'hD5: sbox_out = `SBOX2_ELEMENT_213;
			8'hD6: sbox_out = `SBOX2_ELEMENT_214;
			8'hD7: sbox_out = `SBOX2_ELEMENT_215;
			8'hD8: sbox_out = `SBOX2_ELEMENT_216;
			8'hD9: sbox_out = `SBOX2_ELEMENT_217;
			8'hDA: sbox_out = `SBOX2_ELEMENT_218;
			8'hDB: sbox_out = `SBOX2_ELEMENT_219;
			8'hDC: sbox_out = `SBOX2_ELEMENT_220;
			8'hDD: sbox_out = `SBOX2_ELEMENT_221;
			8'hDE: sbox_out = `SBOX2_ELEMENT_222;
			8'hDF: sbox_out = `SBOX2_ELEMENT_223;
			8'hE0: sbox_out = `SBOX2_ELEMENT_224;
			8'hE1: sbox_out = `SBOX2_ELEMENT_225;
			8'hE2: sbox_out = `SBOX2_ELEMENT_226;
			8'hE3: sbox_out = `SBOX2_ELEMENT_227;
			8'hE4: sbox_out = `SBOX2_ELEMENT_228;
			8'hE5: sbox_out = `SBOX2_ELEMENT_229;
			8'hE6: sbox_out = `SBOX2_ELEMENT_230;
			8'hE7: sbox_out = `SBOX2_ELEMENT_231;
			8'hE8: sbox_out = `SBOX2_ELEMENT_232;
			8'hE9: sbox_out = `SBOX2_ELEMENT_233;
			8'hEA: sbox_out = `SBOX2_ELEMENT_234;
			8'hEB: sbox_out = `SBOX2_ELEMENT_235;
			8'hEC: sbox_out = `SBOX2_ELEMENT_236;
			8'hED: sbox_out = `SBOX2_ELEMENT_237;
			8'hEE: sbox_out = `SBOX2_ELEMENT_238;
			8'hEF: sbox_out = `SBOX2_ELEMENT_239;
			8'hF0: sbox_out = `SBOX2_ELEMENT_240;
			8'hF1: sbox_out = `SBOX2_ELEMENT_241;
			8'hF2: sbox_out = `SBOX2_ELEMENT_242;
			8'hF3: sbox_out = `SBOX2_ELEMENT_243;
			8'hF4: sbox_out = `SBOX2_ELEMENT_244;
			8'hF5: sbox_out = `SBOX2_ELEMENT_245;
			8'hF6: sbox_out = `SBOX2_ELEMENT_246;
			8'hF7: sbox_out = `SBOX2_ELEMENT_247;
			8'hF8: sbox_out = `SBOX2_ELEMENT_248;
			8'hF9: sbox_out = `SBOX2_ELEMENT_249;
			8'hFA: sbox_out = `SBOX2_ELEMENT_250;
			8'hFB: sbox_out = `SBOX2_ELEMENT_251;
			8'hFC: sbox_out = `SBOX2_ELEMENT_252;
			8'hFD: sbox_out = `SBOX2_ELEMENT_253;
			8'hFE: sbox_out = `SBOX2_ELEMENT_254;
			8'hFF: sbox_out = `SBOX2_ELEMENT_255;
			default: sbox_out = 32'h0;
		endcase
	end	
endmodule

`endif
