//-----------------------------------------------------------
// Function: Blowfish-128's S-Boxes
//-----------------------------------------------------------
// Author	: Long Le, Manh Nguyen
// Date  	: Feb-5th, 2025
// Description	: Contains 2 Subtitution Boxes, each has 256 elements 32-bit
//-----------------------------------------------------------

function logic [31:0] blowfish128_sbox1(input [7:0] sbox_in);
	case (sbox_in[7:0])
		8'h00: blowfish128_sbox1[31:0] = 32'hD1310BA6;
		8'h01: blowfish128_sbox1[31:0] = 32'h98DFB5AC;
		8'h02: blowfish128_sbox1[31:0] = 32'h2FFD72DB;
		8'h03: blowfish128_sbox1[31:0] = 32'hD01ADFB7;
		8'h04: blowfish128_sbox1[31:0] = 32'hB8E1AFED;
		8'h05: blowfish128_sbox1[31:0] = 32'h6A267E96;
		8'h06: blowfish128_sbox1[31:0] = 32'hBA7C9045;
		8'h07: blowfish128_sbox1[31:0] = 32'hF12C7F99;
		8'h08: blowfish128_sbox1[31:0] = 32'h24A19947;
		8'h09: blowfish128_sbox1[31:0] = 32'hB3916CF7;
		8'h0A: blowfish128_sbox1[31:0] = 32'h0801F2E2;
		8'h0B: blowfish128_sbox1[31:0] = 32'h858EFC16;
		8'h0C: blowfish128_sbox1[31:0] = 32'h636920D8;
		8'h0D: blowfish128_sbox1[31:0] = 32'h71574E69;
		8'h0E: blowfish128_sbox1[31:0] = 32'hA458FEA3;
		8'h0F: blowfish128_sbox1[31:0] = 32'hF4933D7E;
		8'h10: blowfish128_sbox1[31:0] = 32'h0D95748F;
		8'h11: blowfish128_sbox1[31:0] = 32'h728EB658;
		8'h12: blowfish128_sbox1[31:0] = 32'h718BCD58;
		8'h13: blowfish128_sbox1[31:0] = 32'h82154AEE;
		8'h14: blowfish128_sbox1[31:0] = 32'h7B54A41D;
		8'h15: blowfish128_sbox1[31:0] = 32'hC25A59B5;
		8'h16: blowfish128_sbox1[31:0] = 32'h9C30D539;
		8'h17: blowfish128_sbox1[31:0] = 32'h2AF26013;
		8'h18: blowfish128_sbox1[31:0] = 32'hC5D1B023;
		8'h19: blowfish128_sbox1[31:0] = 32'h286085F0;
		8'h1A: blowfish128_sbox1[31:0] = 32'hCA417918;
		8'h1B: blowfish128_sbox1[31:0] = 32'hB8DB38EF;
		8'h1C: blowfish128_sbox1[31:0] = 32'h8E79DCB0;
		8'h1D: blowfish128_sbox1[31:0] = 32'h603A180E;
		8'h1E: blowfish128_sbox1[31:0] = 32'h6C9E0E8B;
		8'h1F: blowfish128_sbox1[31:0] = 32'hB01E8A3E;
		8'h20: blowfish128_sbox1[31:0] = 32'hD71577C1;
		8'h21: blowfish128_sbox1[31:0] = 32'hBD314B27;
		8'h22: blowfish128_sbox1[31:0] = 32'h78AF2FDA;
		8'h23: blowfish128_sbox1[31:0] = 32'h55605C60;
		8'h24: blowfish128_sbox1[31:0] = 32'hE65525F3;
		8'h25: blowfish128_sbox1[31:0] = 32'hAA55AB94;
		8'h26: blowfish128_sbox1[31:0] = 32'h57489862;
		8'h27: blowfish128_sbox1[31:0] = 32'h63E81440;
		8'h28: blowfish128_sbox1[31:0] = 32'h55CA396A;
		8'h29: blowfish128_sbox1[31:0] = 32'h2AAB10B6;
		8'h2A: blowfish128_sbox1[31:0] = 32'hB4CC5C34;
		8'h2B: blowfish128_sbox1[31:0] = 32'h1141E8CE;
		8'h2C: blowfish128_sbox1[31:0] = 32'hA15486AF;
		8'h2D: blowfish128_sbox1[31:0] = 32'h7C72E993;
		8'h2E: blowfish128_sbox1[31:0] = 32'hB3EE1411;
		8'h2F: blowfish128_sbox1[31:0] = 32'h636FBC2A;
		8'h30: blowfish128_sbox1[31:0] = 32'h2BA9C55D;
		8'h31: blowfish128_sbox1[31:0] = 32'h741831F6;
		8'h32: blowfish128_sbox1[31:0] = 32'hCE5C3E16;
		8'h33: blowfish128_sbox1[31:0] = 32'h9B87931E;
		8'h34: blowfish128_sbox1[31:0] = 32'hAFD6BA33;
		8'h35: blowfish128_sbox1[31:0] = 32'h6C24CF5C;
		8'h36: blowfish128_sbox1[31:0] = 32'h7A325381;
		8'h37: blowfish128_sbox1[31:0] = 32'h28958677;
		8'h38: blowfish128_sbox1[31:0] = 32'h3B8F4898;
		8'h39: blowfish128_sbox1[31:0] = 32'h6B4BB9AF;
		8'h3A: blowfish128_sbox1[31:0] = 32'hC4BFE81B;
		8'h3B: blowfish128_sbox1[31:0] = 32'h66282193;
		8'h3C: blowfish128_sbox1[31:0] = 32'h61D809CC;
		8'h3D: blowfish128_sbox1[31:0] = 32'hFB21A991;
		8'h3E: blowfish128_sbox1[31:0] = 32'h487CAC60;
		8'h3F: blowfish128_sbox1[31:0] = 32'h5DEC8032;
		8'h40: blowfish128_sbox1[31:0] = 32'hEF845D5D;
		8'h41: blowfish128_sbox1[31:0] = 32'hE98575B1;
		8'h42: blowfish128_sbox1[31:0] = 32'hDC262302;
		8'h43: blowfish128_sbox1[31:0] = 32'hEB651B88;
		8'h44: blowfish128_sbox1[31:0] = 32'h23893E81;
		8'h45: blowfish128_sbox1[31:0] = 32'hD396ACC5;
		8'h46: blowfish128_sbox1[31:0] = 32'h0F6D6FF3;
		8'h47: blowfish128_sbox1[31:0] = 32'h83F44239;
		8'h48: blowfish128_sbox1[31:0] = 32'h2E0B4482;
		8'h49: blowfish128_sbox1[31:0] = 32'hA4842004;
		8'h4A: blowfish128_sbox1[31:0] = 32'h69C8F04A;
		8'h4B: blowfish128_sbox1[31:0] = 32'h9E1F9B5E;
		8'h4C: blowfish128_sbox1[31:0] = 32'h21C66842;
		8'h4D: blowfish128_sbox1[31:0] = 32'hF6E96C9A;
		8'h4E: blowfish128_sbox1[31:0] = 32'h670C9C61;
		8'h4F: blowfish128_sbox1[31:0] = 32'hABD388F0;
		8'h50: blowfish128_sbox1[31:0] = 32'h6A51A0D2;
		8'h51: blowfish128_sbox1[31:0] = 32'hD8542F68;
		8'h52: blowfish128_sbox1[31:0] = 32'h960FA728;
		8'h53: blowfish128_sbox1[31:0] = 32'hAB5133A3;
		8'h54: blowfish128_sbox1[31:0] = 32'h6EEF0B6C;
		8'h55: blowfish128_sbox1[31:0] = 32'h137A3BE4;
		8'h56: blowfish128_sbox1[31:0] = 32'hBA3BF050;
		8'h57: blowfish128_sbox1[31:0] = 32'h7EFB2A98;
		8'h58: blowfish128_sbox1[31:0] = 32'hA1F1651D;
		8'h59: blowfish128_sbox1[31:0] = 32'h39AF0176;
		8'h5A: blowfish128_sbox1[31:0] = 32'h66CA593E;
		8'h5B: blowfish128_sbox1[31:0] = 32'h82430E88;
		8'h5C: blowfish128_sbox1[31:0] = 32'h8CEE8619;
		8'h5D: blowfish128_sbox1[31:0] = 32'h456F9FB4;
		8'h5E: blowfish128_sbox1[31:0] = 32'h7D84A5C3;
		8'h5F: blowfish128_sbox1[31:0] = 32'h3B8B5EBE;
		8'h60: blowfish128_sbox1[31:0] = 32'hE06F75D8;
		8'h61: blowfish128_sbox1[31:0] = 32'h85C12073;
		8'h62: blowfish128_sbox1[31:0] = 32'h401A449F;
		8'h63: blowfish128_sbox1[31:0] = 32'h56C16AA6;
		8'h64: blowfish128_sbox1[31:0] = 32'h4ED3AA62;
		8'h65: blowfish128_sbox1[31:0] = 32'h363F7706;
		8'h66: blowfish128_sbox1[31:0] = 32'h1BFEDF72;
		8'h67: blowfish128_sbox1[31:0] = 32'h429B023D;
		8'h68: blowfish128_sbox1[31:0] = 32'h37D0D724;
		8'h69: blowfish128_sbox1[31:0] = 32'hD00A1248;
		8'h6A: blowfish128_sbox1[31:0] = 32'hDB0FEAD3;
		8'h6B: blowfish128_sbox1[31:0] = 32'h49F1C09B;
		8'h6C: blowfish128_sbox1[31:0] = 32'h075372C9;
		8'h6D: blowfish128_sbox1[31:0] = 32'h80991B7B;
		8'h6E: blowfish128_sbox1[31:0] = 32'h25D479D8;
		8'h6F: blowfish128_sbox1[31:0] = 32'hF6E8DEF7;
		8'h70: blowfish128_sbox1[31:0] = 32'hE3FE501A;
		8'h71: blowfish128_sbox1[31:0] = 32'hB6794C3B;
		8'h72: blowfish128_sbox1[31:0] = 32'h976CE0BD;
		8'h73: blowfish128_sbox1[31:0] = 32'h04C006BA;
		8'h74: blowfish128_sbox1[31:0] = 32'hC1A94FB6;
		8'h75: blowfish128_sbox1[31:0] = 32'h409F60C4;
		8'h76: blowfish128_sbox1[31:0] = 32'h5E5C9EC2;
		8'h77: blowfish128_sbox1[31:0] = 32'h196A2463;
		8'h78: blowfish128_sbox1[31:0] = 32'h68FB6FAF;
		8'h79: blowfish128_sbox1[31:0] = 32'h3E6C53B5;
		8'h7A: blowfish128_sbox1[31:0] = 32'h1339B2EB;
		8'h7B: blowfish128_sbox1[31:0] = 32'h3B52EC6F;
		8'h7C: blowfish128_sbox1[31:0] = 32'h6DFC511F;
		8'h7D: blowfish128_sbox1[31:0] = 32'h9B30952C;
		8'h7E: blowfish128_sbox1[31:0] = 32'hCC814544;
		8'h7F: blowfish128_sbox1[31:0] = 32'hAF5EBD09;
		8'h80: blowfish128_sbox1[31:0] = 32'hBEE3D004;
		8'h81: blowfish128_sbox1[31:0] = 32'hDE334AFD;
		8'h82: blowfish128_sbox1[31:0] = 32'h660F2807;
		8'h83: blowfish128_sbox1[31:0] = 32'h192E4BB3;
		8'h84: blowfish128_sbox1[31:0] = 32'hC0CBA857;
		8'h85: blowfish128_sbox1[31:0] = 32'h45C8740F;
		8'h86: blowfish128_sbox1[31:0] = 32'hD20B5F39;
		8'h87: blowfish128_sbox1[31:0] = 32'hB9D3FBDB;
		8'h88: blowfish128_sbox1[31:0] = 32'h5579C0BD;
		8'h89: blowfish128_sbox1[31:0] = 32'h1A60320A;
		8'h8A: blowfish128_sbox1[31:0] = 32'hD6A100C6;
		8'h8B: blowfish128_sbox1[31:0] = 32'h402C7279;
		8'h8C: blowfish128_sbox1[31:0] = 32'h679F25FE;
		8'h8D: blowfish128_sbox1[31:0] = 32'hFB1FA3CC;
		8'h8E: blowfish128_sbox1[31:0] = 32'h8EA5E9F8;
		8'h8F: blowfish128_sbox1[31:0] = 32'hDB3222F8;
		8'h90: blowfish128_sbox1[31:0] = 32'h3C7516DF;
		8'h91: blowfish128_sbox1[31:0] = 32'hFD616B15;
		8'h92: blowfish128_sbox1[31:0] = 32'h2F501EC8;
		8'h93: blowfish128_sbox1[31:0] = 32'hAD0552AB;
		8'h94: blowfish128_sbox1[31:0] = 32'h323DB5FA;
		8'h95: blowfish128_sbox1[31:0] = 32'hFD238760;
		8'h96: blowfish128_sbox1[31:0] = 32'h53317B48;
		8'h97: blowfish128_sbox1[31:0] = 32'h3E00DF82;
		8'h98: blowfish128_sbox1[31:0] = 32'h9E5C57BB;
		8'h99: blowfish128_sbox1[31:0] = 32'hCA6F8CA0;
		8'h9A: blowfish128_sbox1[31:0] = 32'h1A87562E;
		8'h9B: blowfish128_sbox1[31:0] = 32'hDF1769DB;
		8'h9C: blowfish128_sbox1[31:0] = 32'hD542A8F6;
		8'h9D: blowfish128_sbox1[31:0] = 32'h287EFFC3;
		8'h9E: blowfish128_sbox1[31:0] = 32'hAC6732C6;
		8'h9F: blowfish128_sbox1[31:0] = 32'h8C4F5573;
		8'hA0: blowfish128_sbox1[31:0] = 32'h695B27B0;
		8'hA1: blowfish128_sbox1[31:0] = 32'hBBCA58C8;
		8'hA2: blowfish128_sbox1[31:0] = 32'hE1FFA35D;
		8'hA3: blowfish128_sbox1[31:0] = 32'hB8F011A0;
		8'hA4: blowfish128_sbox1[31:0] = 32'h10FA3D98;
		8'hA5: blowfish128_sbox1[31:0] = 32'hFD2183B8;
		8'hA6: blowfish128_sbox1[31:0] = 32'h4AFCB56C;
		8'hA7: blowfish128_sbox1[31:0] = 32'h2DD1D35B;
		8'hA8: blowfish128_sbox1[31:0] = 32'h9A53E479;
		8'hA9: blowfish128_sbox1[31:0] = 32'hB6F84565;
		8'hAA: blowfish128_sbox1[31:0] = 32'hD28E49BC;
		8'hAB: blowfish128_sbox1[31:0] = 32'h4BFB9790;
		8'hAC: blowfish128_sbox1[31:0] = 32'hE1DDF2DA;
		8'hAD: blowfish128_sbox1[31:0] = 32'hA4CB7E33;
		8'hAE: blowfish128_sbox1[31:0] = 32'h62FB1341;
		8'hAF: blowfish128_sbox1[31:0] = 32'hCEE4C6E8;
		8'hB0: blowfish128_sbox1[31:0] = 32'hEF20CADA;
		8'hB1: blowfish128_sbox1[31:0] = 32'h36774C01;
		8'hB2: blowfish128_sbox1[31:0] = 32'hD07E9EFE;
		8'hB3: blowfish128_sbox1[31:0] = 32'h2BF11FB4;
		8'hB4: blowfish128_sbox1[31:0] = 32'h95DBDA4D;
		8'hB5: blowfish128_sbox1[31:0] = 32'hAE909198;
		8'hB6: blowfish128_sbox1[31:0] = 32'hEAAD8E71;
		8'hB7: blowfish128_sbox1[31:0] = 32'h6B93D5A0;
		8'hB8: blowfish128_sbox1[31:0] = 32'hD08ED1D0;
		8'hB9: blowfish128_sbox1[31:0] = 32'hAFC725E0;
		8'hBA: blowfish128_sbox1[31:0] = 32'h8E3C5B2F;
		8'hBB: blowfish128_sbox1[31:0] = 32'h8E7594B7;
		8'hBC: blowfish128_sbox1[31:0] = 32'h8FF6E2FB;
		8'hBD: blowfish128_sbox1[31:0] = 32'hF2122B64;
		8'hBE: blowfish128_sbox1[31:0] = 32'h8888B812;
		8'hBF: blowfish128_sbox1[31:0] = 32'h900DF01C;
		8'hC0: blowfish128_sbox1[31:0] = 32'h4FAD5EA0;
		8'hC1: blowfish128_sbox1[31:0] = 32'h688FC31C;
		8'hC2: blowfish128_sbox1[31:0] = 32'hD1CFF191;
		8'hC3: blowfish128_sbox1[31:0] = 32'hB3A8C1AD;
		8'hC4: blowfish128_sbox1[31:0] = 32'h2F2F2218;
		8'hC5: blowfish128_sbox1[31:0] = 32'hBE0E1777;
		8'hC6: blowfish128_sbox1[31:0] = 32'hEA752DFE;
		8'hC7: blowfish128_sbox1[31:0] = 32'h8B021FA1;
		8'hC8: blowfish128_sbox1[31:0] = 32'hE5A0CC0F;
		8'hC9: blowfish128_sbox1[31:0] = 32'hB56F74E8;
		8'hCA: blowfish128_sbox1[31:0] = 32'h18ACF3D6;
		8'hCB: blowfish128_sbox1[31:0] = 32'hCE89E299;
		8'hCC: blowfish128_sbox1[31:0] = 32'hB4A84FE0;
		8'hCD: blowfish128_sbox1[31:0] = 32'hFD13E0B7;
		8'hCE: blowfish128_sbox1[31:0] = 32'h7CC43B81;
		8'hCF: blowfish128_sbox1[31:0] = 32'hD2ADA8D9;
		8'hD0: blowfish128_sbox1[31:0] = 32'h165FA266;
		8'hD1: blowfish128_sbox1[31:0] = 32'h80957705;
		8'hD2: blowfish128_sbox1[31:0] = 32'h93CC7314;
		8'hD3: blowfish128_sbox1[31:0] = 32'h211A1477;
		8'hD4: blowfish128_sbox1[31:0] = 32'hE6AD2065;
		8'hD5: blowfish128_sbox1[31:0] = 32'h77B5FA86;
		8'hD6: blowfish128_sbox1[31:0] = 32'hC75442F5;
		8'hD7: blowfish128_sbox1[31:0] = 32'hFB9D35CF;
		8'hD8: blowfish128_sbox1[31:0] = 32'hEBCDAF0C;
		8'hD9: blowfish128_sbox1[31:0] = 32'h7B3E89A0;
		8'hDA: blowfish128_sbox1[31:0] = 32'hD6411BD3;
		8'hDB: blowfish128_sbox1[31:0] = 32'hAE1E7E49;
		8'hDC: blowfish128_sbox1[31:0] = 32'h00250E2D;
		8'hDD: blowfish128_sbox1[31:0] = 32'h2071B35E;
		8'hDE: blowfish128_sbox1[31:0] = 32'h226800BB;
		8'hDF: blowfish128_sbox1[31:0] = 32'h57B8E0AF;
		8'hE0: blowfish128_sbox1[31:0] = 32'h2464369B;
		8'hE1: blowfish128_sbox1[31:0] = 32'hF009B91E;
		8'hE2: blowfish128_sbox1[31:0] = 32'h5563911D;
		8'hE3: blowfish128_sbox1[31:0] = 32'h59DFA6AA;
		8'hE4: blowfish128_sbox1[31:0] = 32'h78C14389;
		8'hE5: blowfish128_sbox1[31:0] = 32'hD95A537F;
		8'hE6: blowfish128_sbox1[31:0] = 32'h207D5BA2;
		8'hE7: blowfish128_sbox1[31:0] = 32'h02E5B9C5;
		8'hE8: blowfish128_sbox1[31:0] = 32'h83260376;
		8'hE9: blowfish128_sbox1[31:0] = 32'h6295CFA9;
		8'hEA: blowfish128_sbox1[31:0] = 32'h11C81968;
		8'hEB: blowfish128_sbox1[31:0] = 32'h4E734A41;
		8'hEC: blowfish128_sbox1[31:0] = 32'hB3472DCA;
		8'hED: blowfish128_sbox1[31:0] = 32'h7B14A94A;
		8'hEE: blowfish128_sbox1[31:0] = 32'h1B510052;
		8'hEF: blowfish128_sbox1[31:0] = 32'h9A532915;
		8'hF0: blowfish128_sbox1[31:0] = 32'hD60F573F;
		8'hF1: blowfish128_sbox1[31:0] = 32'hBC9BC6E4;
		8'hF2: blowfish128_sbox1[31:0] = 32'h2B60A476;
		8'hF3: blowfish128_sbox1[31:0] = 32'h81E67400;
		8'hF4: blowfish128_sbox1[31:0] = 32'h08BA6FB5;
		8'hF5: blowfish128_sbox1[31:0] = 32'h571BE91F;
		8'hF6: blowfish128_sbox1[31:0] = 32'hF296EC6B;
		8'hF7: blowfish128_sbox1[31:0] = 32'h2A0DD915;
		8'hF8: blowfish128_sbox1[31:0] = 32'hB6636521;
		8'hF9: blowfish128_sbox1[31:0] = 32'hE7B9F9B6;
		8'hFA: blowfish128_sbox1[31:0] = 32'hFF34052E;
		8'hFB: blowfish128_sbox1[31:0] = 32'hC5855664;
		8'hFC: blowfish128_sbox1[31:0] = 32'h53B02D5D;
		8'hFD: blowfish128_sbox1[31:0] = 32'hA99F8FA1;
		8'hFE: blowfish128_sbox1[31:0] = 32'h08BA4799;
		8'hFF: blowfish128_sbox1[31:0] = 32'h6E85076A;
		default: blowfish128_sbox1[31:0] = 32'hXXXXXXXX;
	endcase
endfunction: blowfish128_sbox1

function logic [31:0] blowfish128_sbox2(input [7:0] sbox_in);
	case(sbox_in[7:0])
		8'h00: blowfish128_sbox2[31:0] = 32'h4B7A70E9;
		8'h01: blowfish128_sbox2[31:0] = 32'hB5B32944;
		8'h02: blowfish128_sbox2[31:0] = 32'hDB75092E;
		8'h03: blowfish128_sbox2[31:0] = 32'hC4192623;
		8'h04: blowfish128_sbox2[31:0] = 32'hAD6EA6B0;
		8'h05: blowfish128_sbox2[31:0] = 32'h49A7DF7D;
		8'h06: blowfish128_sbox2[31:0] = 32'h9CEE60B8;
		8'h07: blowfish128_sbox2[31:0] = 32'h8FEDB266;
		8'h08: blowfish128_sbox2[31:0] = 32'hECAA8C71;
		8'h09: blowfish128_sbox2[31:0] = 32'h699A17FF;
		8'h0A: blowfish128_sbox2[31:0] = 32'h5664526C;
		8'h0B: blowfish128_sbox2[31:0] = 32'hC2B19EE1;
		8'h0C: blowfish128_sbox2[31:0] = 32'h193602A5;
		8'h0D: blowfish128_sbox2[31:0] = 32'h75094C29;
		8'h0E: blowfish128_sbox2[31:0] = 32'hA0591340;
		8'h0F: blowfish128_sbox2[31:0] = 32'hE4183A3E;
		8'h10: blowfish128_sbox2[31:0] = 32'h3F54989A;
		8'h11: blowfish128_sbox2[31:0] = 32'h5B429D65;
		8'h12: blowfish128_sbox2[31:0] = 32'h6B8FE4D6;
		8'h13: blowfish128_sbox2[31:0] = 32'h99F73FD6;
		8'h14: blowfish128_sbox2[31:0] = 32'hA1D29C07;
		8'h15: blowfish128_sbox2[31:0] = 32'hEFE830F5;
		8'h16: blowfish128_sbox2[31:0] = 32'h4D2D38E6;
		8'h17: blowfish128_sbox2[31:0] = 32'hF0255DC1;
		8'h18: blowfish128_sbox2[31:0] = 32'h4CDD2086;
		8'h19: blowfish128_sbox2[31:0] = 32'h8470EB26;
		8'h1A: blowfish128_sbox2[31:0] = 32'h6382E9C6;
		8'h1B: blowfish128_sbox2[31:0] = 32'h021ECC5E;
		8'h1C: blowfish128_sbox2[31:0] = 32'h09686B3F;
		8'h1D: blowfish128_sbox2[31:0] = 32'h3EBAEFC9;
		8'h1E: blowfish128_sbox2[31:0] = 32'h3C971814;
		8'h1F: blowfish128_sbox2[31:0] = 32'h6B6A70A1;
		8'h20: blowfish128_sbox2[31:0] = 32'h687F3584;
		8'h21: blowfish128_sbox2[31:0] = 32'h52A0E286;
		8'h22: blowfish128_sbox2[31:0] = 32'hB79C5305;
		8'h23: blowfish128_sbox2[31:0] = 32'hAA500737;
		8'h24: blowfish128_sbox2[31:0] = 32'h3E07841C;
		8'h25: blowfish128_sbox2[31:0] = 32'h7FDEAE5C;
		8'h26: blowfish128_sbox2[31:0] = 32'h8E7D44EC;
		8'h27: blowfish128_sbox2[31:0] = 32'h5716F2B8;
		8'h28: blowfish128_sbox2[31:0] = 32'hB03ADA37;
		8'h29: blowfish128_sbox2[31:0] = 32'hF0500C0D;
		8'h2A: blowfish128_sbox2[31:0] = 32'hF01C1F04;
		8'h2B: blowfish128_sbox2[31:0] = 32'h0200B3FF;
		8'h2C: blowfish128_sbox2[31:0] = 32'hAE0CF51A;
		8'h2D: blowfish128_sbox2[31:0] = 32'h3CB574B2;
		8'h2E: blowfish128_sbox2[31:0] = 32'h25837A58;
		8'h2F: blowfish128_sbox2[31:0] = 32'hDC0921BD;
		8'h30: blowfish128_sbox2[31:0] = 32'hD19113F9;
		8'h31: blowfish128_sbox2[31:0] = 32'h7CA92FF6;
		8'h32: blowfish128_sbox2[31:0] = 32'h94324773;
		8'h33: blowfish128_sbox2[31:0] = 32'h22F54701;
		8'h34: blowfish128_sbox2[31:0] = 32'h3AE5E581;
		8'h35: blowfish128_sbox2[31:0] = 32'h37C2DADC;
		8'h36: blowfish128_sbox2[31:0] = 32'hC8B57634;
		8'h37: blowfish128_sbox2[31:0] = 32'h9AF3DDA7;
		8'h38: blowfish128_sbox2[31:0] = 32'hA9446146;
		8'h39: blowfish128_sbox2[31:0] = 32'h0FD0030E;
		8'h3A: blowfish128_sbox2[31:0] = 32'hECC8C73E;
		8'h3B: blowfish128_sbox2[31:0] = 32'hA4751E41;
		8'h3C: blowfish128_sbox2[31:0] = 32'hE238CD99;
		8'h3D: blowfish128_sbox2[31:0] = 32'h3BEA0E2F;
		8'h3E: blowfish128_sbox2[31:0] = 32'h3280BBA1;
		8'h3F: blowfish128_sbox2[31:0] = 32'h183EB331;
		8'h40: blowfish128_sbox2[31:0] = 32'h4E548B38;
		8'h41: blowfish128_sbox2[31:0] = 32'h4F6DB908;
		8'h42: blowfish128_sbox2[31:0] = 32'h6F420D03;
		8'h43: blowfish128_sbox2[31:0] = 32'hF60A04BF;
		8'h44: blowfish128_sbox2[31:0] = 32'h2CB81290;
		8'h45: blowfish128_sbox2[31:0] = 32'h24977C79;
		8'h46: blowfish128_sbox2[31:0] = 32'h5679B072;
		8'h47: blowfish128_sbox2[31:0] = 32'hBCAF89AF;
		8'h48: blowfish128_sbox2[31:0] = 32'hDE9A771F;
		8'h49: blowfish128_sbox2[31:0] = 32'hD9930810;
		8'h4A: blowfish128_sbox2[31:0] = 32'hB38BAE12;
		8'h4B: blowfish128_sbox2[31:0] = 32'hDCCF3F2E;
		8'h4C: blowfish128_sbox2[31:0] = 32'h5512721F;
		8'h4D: blowfish128_sbox2[31:0] = 32'h2E6B7124;
		8'h4E: blowfish128_sbox2[31:0] = 32'h501ADDE6;
		8'h4F: blowfish128_sbox2[31:0] = 32'h9F84CD87;
		8'h50: blowfish128_sbox2[31:0] = 32'h7A584718;
		8'h51: blowfish128_sbox2[31:0] = 32'h7408DA17;
		8'h52: blowfish128_sbox2[31:0] = 32'hBC9F9ABC;
		8'h53: blowfish128_sbox2[31:0] = 32'hE94B7D8C;
		8'h54: blowfish128_sbox2[31:0] = 32'hEC7AEC3A;
		8'h55: blowfish128_sbox2[31:0] = 32'hDB851DFA;
		8'h56: blowfish128_sbox2[31:0] = 32'h63094366;
		8'h57: blowfish128_sbox2[31:0] = 32'hC464C3D2;
		8'h58: blowfish128_sbox2[31:0] = 32'hEF1C1847;
		8'h59: blowfish128_sbox2[31:0] = 32'h3215D908;
		8'h5A: blowfish128_sbox2[31:0] = 32'hDD433B37;
		8'h5B: blowfish128_sbox2[31:0] = 32'h24C2BA16;
		8'h5C: blowfish128_sbox2[31:0] = 32'h12A14D43;
		8'h5D: blowfish128_sbox2[31:0] = 32'h2A65C451;
		8'h5E: blowfish128_sbox2[31:0] = 32'h50940002;
		8'h5F: blowfish128_sbox2[31:0] = 32'h133AE4DD;
		8'h60: blowfish128_sbox2[31:0] = 32'h71DFF89E;
		8'h61: blowfish128_sbox2[31:0] = 32'h10314E55;
		8'h62: blowfish128_sbox2[31:0] = 32'h81AC77D6;
		8'h63: blowfish128_sbox2[31:0] = 32'h5F11199B;
		8'h64: blowfish128_sbox2[31:0] = 32'h043556F1;
		8'h65: blowfish128_sbox2[31:0] = 32'hD7A3C76B;
		8'h66: blowfish128_sbox2[31:0] = 32'h3C11183B;
		8'h67: blowfish128_sbox2[31:0] = 32'h5924A509;
		8'h68: blowfish128_sbox2[31:0] = 32'hF28FE6ED;
		8'h69: blowfish128_sbox2[31:0] = 32'h97F1FBFA;
		8'h6A: blowfish128_sbox2[31:0] = 32'h9EBABF2C;
		8'h6B: blowfish128_sbox2[31:0] = 32'h1E153C6E;
		8'h6C: blowfish128_sbox2[31:0] = 32'h86E34570;
		8'h6D: blowfish128_sbox2[31:0] = 32'hEAE96FB1;
		8'h6E: blowfish128_sbox2[31:0] = 32'h860E5E0A;
		8'h6F: blowfish128_sbox2[31:0] = 32'h5A3E2AB3;
		8'h70: blowfish128_sbox2[31:0] = 32'h771FE71C;
		8'h71: blowfish128_sbox2[31:0] = 32'h4E3D06FA;
		8'h72: blowfish128_sbox2[31:0] = 32'h2965DCB9;
		8'h73: blowfish128_sbox2[31:0] = 32'h99E71D0F;
		8'h74: blowfish128_sbox2[31:0] = 32'h803E89D6;
		8'h75: blowfish128_sbox2[31:0] = 32'h5266C825;
		8'h76: blowfish128_sbox2[31:0] = 32'h2E4CC978;
		8'h77: blowfish128_sbox2[31:0] = 32'h9C10B36A;
		8'h78: blowfish128_sbox2[31:0] = 32'hC6150EBA;
		8'h79: blowfish128_sbox2[31:0] = 32'h94E2EA78;
		8'h7A: blowfish128_sbox2[31:0] = 32'hA5FC3C53;
		8'h7B: blowfish128_sbox2[31:0] = 32'h1E0A2DF4;
		8'h7C: blowfish128_sbox2[31:0] = 32'hF2F74EA7;
		8'h7D: blowfish128_sbox2[31:0] = 32'h361D2B3D;
		8'h7E: blowfish128_sbox2[31:0] = 32'h1939260F;
		8'h7F: blowfish128_sbox2[31:0] = 32'h19C27960;
		8'h80: blowfish128_sbox2[31:0] = 32'h5223A708;
		8'h81: blowfish128_sbox2[31:0] = 32'hF71312B6;
		8'h82: blowfish128_sbox2[31:0] = 32'hEBADFE6E;
		8'h83: blowfish128_sbox2[31:0] = 32'hEAC31F66;
		8'h84: blowfish128_sbox2[31:0] = 32'hE3BC4595;
		8'h85: blowfish128_sbox2[31:0] = 32'hA67BC883;
		8'h86: blowfish128_sbox2[31:0] = 32'hB17F37D1;
		8'h87: blowfish128_sbox2[31:0] = 32'h018CFF28;
		8'h88: blowfish128_sbox2[31:0] = 32'hC332DDEF;
		8'h89: blowfish128_sbox2[31:0] = 32'hBE6C5AA5;
		8'h8A: blowfish128_sbox2[31:0] = 32'h65582185;
		8'h8B: blowfish128_sbox2[31:0] = 32'h68AB9802;
		8'h8C: blowfish128_sbox2[31:0] = 32'hEECEA50F;
		8'h8D: blowfish128_sbox2[31:0] = 32'hDB2F953B;
		8'h8E: blowfish128_sbox2[31:0] = 32'h2AEF7DAD;
		8'h8F: blowfish128_sbox2[31:0] = 32'h5B6E2F84;
		8'h90: blowfish128_sbox2[31:0] = 32'h1521B628;
		8'h91: blowfish128_sbox2[31:0] = 32'h29076170;
		8'h92: blowfish128_sbox2[31:0] = 32'hECDD4775;
		8'h93: blowfish128_sbox2[31:0] = 32'h619F1510;
		8'h94: blowfish128_sbox2[31:0] = 32'h13CCA830;
		8'h95: blowfish128_sbox2[31:0] = 32'hEB61BD96;
		8'h96: blowfish128_sbox2[31:0] = 32'h0334FE1E;
		8'h97: blowfish128_sbox2[31:0] = 32'hAA0363CF;
		8'h98: blowfish128_sbox2[31:0] = 32'hB5735C90;
		8'h99: blowfish128_sbox2[31:0] = 32'h4C70A239;
		8'h9A: blowfish128_sbox2[31:0] = 32'hD59E9E0B;
		8'h9B: blowfish128_sbox2[31:0] = 32'hCBAADE14;
		8'h9C: blowfish128_sbox2[31:0] = 32'hEECC86BC;
		8'h9D: blowfish128_sbox2[31:0] = 32'h60622CA7;
		8'h9E: blowfish128_sbox2[31:0] = 32'h9CAB5CAB;
		8'h9F: blowfish128_sbox2[31:0] = 32'hB2F3846E;
		8'hA0: blowfish128_sbox2[31:0] = 32'h648B1EAF;
		8'hA1: blowfish128_sbox2[31:0] = 32'h19BDF0CA;
		8'hA2: blowfish128_sbox2[31:0] = 32'hA02369B9;
		8'hA3: blowfish128_sbox2[31:0] = 32'h655ABB50;
		8'hA4: blowfish128_sbox2[31:0] = 32'h40685A32;
		8'hA5: blowfish128_sbox2[31:0] = 32'h3C2AB4B3;
		8'hA6: blowfish128_sbox2[31:0] = 32'h319EE9D5;
		8'hA7: blowfish128_sbox2[31:0] = 32'hC021B8F7;
		8'hA8: blowfish128_sbox2[31:0] = 32'h9B540B19;
		8'hA9: blowfish128_sbox2[31:0] = 32'h875FA099;
		8'hAA: blowfish128_sbox2[31:0] = 32'h95F7997E;
		8'hAB: blowfish128_sbox2[31:0] = 32'h623D7DA8;
		8'hAC: blowfish128_sbox2[31:0] = 32'hF837889A;
		8'hAD: blowfish128_sbox2[31:0] = 32'h97E32D77;
		8'hAE: blowfish128_sbox2[31:0] = 32'h11ED935F;
		8'hAF: blowfish128_sbox2[31:0] = 32'h16681281;
		8'hB0: blowfish128_sbox2[31:0] = 32'h0E358829;
		8'hB1: blowfish128_sbox2[31:0] = 32'hC7E61FD6;
		8'hB2: blowfish128_sbox2[31:0] = 32'h96DEDFA1;
		8'hB3: blowfish128_sbox2[31:0] = 32'h7858BA99;
		8'hB4: blowfish128_sbox2[31:0] = 32'h57F584A5;
		8'hB5: blowfish128_sbox2[31:0] = 32'h1B227263;
		8'hB6: blowfish128_sbox2[31:0] = 32'h9B83C3FF;
		8'hB7: blowfish128_sbox2[31:0] = 32'h1AC24696;
		8'hB8: blowfish128_sbox2[31:0] = 32'hCDB30AEB;
		8'hB9: blowfish128_sbox2[31:0] = 32'h532E3054;
		8'hBA: blowfish128_sbox2[31:0] = 32'h8FD948E4;
		8'hBB: blowfish128_sbox2[31:0] = 32'h6DBC3128;
		8'hBC: blowfish128_sbox2[31:0] = 32'h58EBF2EF;
		8'hBD: blowfish128_sbox2[31:0] = 32'h34C6FFEA;
		8'hBE: blowfish128_sbox2[31:0] = 32'hFE28ED61;
		8'hBF: blowfish128_sbox2[31:0] = 32'hEE7C3C73;
		8'hC0: blowfish128_sbox2[31:0] = 32'h5D4A14D9;
		8'hC1: blowfish128_sbox2[31:0] = 32'hE864B7E3;
		8'hC2: blowfish128_sbox2[31:0] = 32'h42105D14;
		8'hC3: blowfish128_sbox2[31:0] = 32'h203E13E0;
		8'hC4: blowfish128_sbox2[31:0] = 32'h45EEE2B6;
		8'hC5: blowfish128_sbox2[31:0] = 32'hA3AAABEA;
		8'hC6: blowfish128_sbox2[31:0] = 32'hDB6C4F15;
		8'hC7: blowfish128_sbox2[31:0] = 32'hFACB4FD0;
		8'hC8: blowfish128_sbox2[31:0] = 32'hC742F442;
		8'hC9: blowfish128_sbox2[31:0] = 32'hEF6ABBB5;
		8'hCA: blowfish128_sbox2[31:0] = 32'h654F3B1D;
		8'hCB: blowfish128_sbox2[31:0] = 32'h41CD2105;
		8'hCC: blowfish128_sbox2[31:0] = 32'hD81E799E;
		8'hCD: blowfish128_sbox2[31:0] = 32'h86854DC7;
		8'hCE: blowfish128_sbox2[31:0] = 32'hE44B476A;
		8'hCF: blowfish128_sbox2[31:0] = 32'h3D816250;
		8'hD0: blowfish128_sbox2[31:0] = 32'hCF62A1F2;
		8'hD1: blowfish128_sbox2[31:0] = 32'h5B8D2646;
		8'hD2: blowfish128_sbox2[31:0] = 32'hFC8883A0;
		8'hD3: blowfish128_sbox2[31:0] = 32'hC1C7B6A3;
		8'hD4: blowfish128_sbox2[31:0] = 32'h7F1524C3;
		8'hD5: blowfish128_sbox2[31:0] = 32'h69CB7492;
		8'hD6: blowfish128_sbox2[31:0] = 32'h47848A0B;
		8'hD7: blowfish128_sbox2[31:0] = 32'h5692B285;
		8'hD8: blowfish128_sbox2[31:0] = 32'h095BBF00;
		8'hD9: blowfish128_sbox2[31:0] = 32'hAD19489D;
		8'hDA: blowfish128_sbox2[31:0] = 32'h1462B174;
		8'hDB: blowfish128_sbox2[31:0] = 32'h23820E00;
		8'hDC: blowfish128_sbox2[31:0] = 32'h58428D2A;
		8'hDD: blowfish128_sbox2[31:0] = 32'h0C55F5EA;
		8'hDE: blowfish128_sbox2[31:0] = 32'h1DADF43E;
		8'hDF: blowfish128_sbox2[31:0] = 32'h233F7061;
		8'hE0: blowfish128_sbox2[31:0] = 32'h3372F092;
		8'hE1: blowfish128_sbox2[31:0] = 32'h8D937E41;
		8'hE2: blowfish128_sbox2[31:0] = 32'hD65FECF1;
		8'hE3: blowfish128_sbox2[31:0] = 32'h6C223BDB;
		8'hE4: blowfish128_sbox2[31:0] = 32'h7CDE3759;
		8'hE5: blowfish128_sbox2[31:0] = 32'hCBEE7460;
		8'hE6: blowfish128_sbox2[31:0] = 32'h4085F2A7;
		8'hE7: blowfish128_sbox2[31:0] = 32'hCE77326E;
		8'hE8: blowfish128_sbox2[31:0] = 32'hA6078084;
		8'hE9: blowfish128_sbox2[31:0] = 32'h19F8509E;
		8'hEA: blowfish128_sbox2[31:0] = 32'hE8EFD855;
		8'hEB: blowfish128_sbox2[31:0] = 32'h61D99735;
		8'hEC: blowfish128_sbox2[31:0] = 32'hA969A7AA;
		8'hED: blowfish128_sbox2[31:0] = 32'hC50C06C2;
		8'hEE: blowfish128_sbox2[31:0] = 32'h5A04ABFC;
		8'hEF: blowfish128_sbox2[31:0] = 32'h800BCADC;
		8'hF0: blowfish128_sbox2[31:0] = 32'h9E447A2E;
		8'hF1: blowfish128_sbox2[31:0] = 32'hC3453484;
		8'hF2: blowfish128_sbox2[31:0] = 32'hFDD56705;
		8'hF3: blowfish128_sbox2[31:0] = 32'h0E1E9EC9;
		8'hF4: blowfish128_sbox2[31:0] = 32'hDB73DBD3;
		8'hF5: blowfish128_sbox2[31:0] = 32'h105588CD;
		8'hF6: blowfish128_sbox2[31:0] = 32'h675FDA79;
		8'hF7: blowfish128_sbox2[31:0] = 32'hE3674340;
		8'hF8: blowfish128_sbox2[31:0] = 32'hC5C43465;
		8'hF9: blowfish128_sbox2[31:0] = 32'h713E38D8;
		8'hFA: blowfish128_sbox2[31:0] = 32'h3D28F89E;
		8'hFB: blowfish128_sbox2[31:0] = 32'hF16DFF20;
		8'hFC: blowfish128_sbox2[31:0] = 32'h153E21E7;
		8'hFD: blowfish128_sbox2[31:0] = 32'h8FB03D4A;
		8'hFE: blowfish128_sbox2[31:0] = 32'hE6E39F2B;
		8'hFF: blowfish128_sbox2[31:0] = 32'hDB83ADF7;
		default: blowfish128_sbox2[31:0] = 32'hXXXXXXXX;
	endcase
endfunction: blowfish128_sbox2
