interface IBR128_if;
	logic Clk;
	logic RstN;
	logic CS;
	logic Write;
	logic Read;
	logic [4:0] Addr;
	logic [31:0] WData;
	logic [31:0] RData;
endinterface
